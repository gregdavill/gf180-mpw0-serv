* NGSPICE file created from serv_0.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_ip_sram__sram256x8m8wm1 abstract view
.subckt gf180mcu_fd_ip_sram__sram256x8m8wm1 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7]
+ CEN CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] GWEN Q[0] Q[1] Q[2] Q[3] Q[4] Q[5]
+ Q[6] Q[7] WEN[0] WEN[1] WEN[2] WEN[3] WEN[4] WEN[5] WEN[6] WEN[7] VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

.subckt serv_0 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_45_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3155_ _0149_ net97 u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2106_ _1282_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout56_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3086_ _0083_ net57 u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _0225_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.raddr\[0\] u_cpu.rf_ram_if.rcnt\[2\]
+ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_39_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2254__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2939_ _0982_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2954__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2621__C _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1693__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2642__B1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2945__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[34\] u_arbiter.i_wb_cpu_rdt\[31\] net145 u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ net27 u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2173__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[68\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1684__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2773__I _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2484__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2236__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1739__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _0845_
+ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2655_ _0560_ _0630_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1606_ _1083_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2586_ _0414_ _0554_ _0739_ _0528_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout127 net130 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1852__I u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout138 net142 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout105 net110 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3207_ _0200_ net54 u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3138_ _0135_ net118 u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1801__B _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3069_ _0066_ net116 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1666__A1 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2091__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3028__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3178__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[2\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ _0511_ _0593_ _0605_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2371_ _0437_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2854__B1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout19_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _0836_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2385__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2638_ u_cpu.cpu.immdec.imm19_12_20\[6\] _0514_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2569_ u_cpu.cpu.immdec.imm30_25\[5\] _0678_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1648__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2845__B1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1639__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2687__I0 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2300__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1940_ _1076_ _1361_ _1364_ u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_124_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1871_ _1248_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1811__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2423_ _0579_ _0590_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2354_ _0501_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2285_ _0415_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2530__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2046__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3216__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2070_ _1246_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2982__S _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2972_ _1011_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1923_ _1347_ _1341_ _1353_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1854_ _1049_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1785_ _1225_ _1229_ u_arbiter.i_wb_cpu_dbus_we _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2406_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2899__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout86_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2337_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2268_ _0438_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2276__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2199_ u_arbiter.i_wb_cpu_rdt\[19\] _0386_ _0355_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2028__A1 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__C _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3239__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2534__C _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[64\] u_scanchain_local.module_data_in\[63\] net147 u_arbiter.o_wb_cpu_adr\[26\]
+ net30 u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _1045_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3240_ u_cpu.cpu.o_wen1 net56 u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3171_ _0165_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2776__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _1321_ net35 _0317_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2053_ _0273_ _0233_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _1250_ _0277_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1906_ _1226_ u_cpu.rf_ram.rdata\[5\] _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2886_ _0474_ _0657_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1837_ _1212_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2981__A2 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1768_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1699_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _1157_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2249__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2421__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1775__A3 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput7 net7 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2488__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2660__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ _0854_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout136_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2671_ _0553_ _0620_ _0710_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1622_ _1095_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3223_ u_cpu.rf_ram_if.wdata0_r\[6\] net45 u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2479__A1 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3154_ _0148_ net100 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2105_ _1213_ _0312_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3085_ _0082_ net57 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_36_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2455__B _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2036_ _0255_ _0258_ _0260_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout49_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3084__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2938_ _1372_ _1377_ _0987_ _1077_ _1063_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2403__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2954__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2869_ _0594_ _0937_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1765__I0 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__B2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2642__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[27\] u_arbiter.i_wb_cpu_rdt\[24\] net143 u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ net28 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_46_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2881__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2633__B2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2633__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2723_ _0826_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2654_ _0709_ _0764_ _0798_ _0799_ _0630_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2585_ _0735_ _0432_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1605_ _1068_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout117 net121 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout106 net110 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout139 net141 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_45_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[12\]_SE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3206_ _0199_ net70 u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3137_ _0134_ net119 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3068_ _0065_ net115 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2019_ _0225_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[2\] _0248_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2624__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[23\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[38\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1666__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2615__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1953__I _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[35\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2370_ _0494_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2985__S _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2854__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2854__B2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3122__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _0833_
+ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2637_ _0484_ _0775_ _0784_ _0653_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2568_ _0511_ _0718_ _0722_ _0514_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1896__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2499_ _0502_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2845__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2073__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1584__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1773__I u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1887__A2 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2533__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2687__I1 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3145__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1948__I _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1870_ _1311_ u_cpu.cpu.ctrl.i_iscomp _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2422_ _0580_ _0581_ _0586_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ _0489_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2284_ _0227_ u_arbiter.i_wb_cpu_rdt\[8\] _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_42_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1999_ net8 _1086_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3018__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1869__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[1\]_CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1768__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2373__B _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2599__I _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2506__B1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2285__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2971_ _1333_ _1335_ u_cpu.rf_ram.rdata\[7\] _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_91_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ u_cpu.rf_ram_if.rdata0\[5\] _1350_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1853_ _1295_ u_cpu.cpu.alu.add_cy_r _1231_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1784_ u_cpu.rf_ram_if.rtrig1 _1227_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_89_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout8 u_arbiter.i_wb_cpu_ack net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2302__I _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _0451_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout79_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1720__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2336_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2267_ _0429_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _0357_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2520__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2276__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2413__S _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3000__I1 u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1711__A1 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2368__B _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2882__I u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2267__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[57\] u_scanchain_local.module_data_in\[56\] net139 u_arbiter.o_wb_cpu_adr\[19\]
+ net23 u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1961__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3170_ _0164_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _0317_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2993__S _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2052_ _1218_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2954_ u_cpu.cpu.decode.co_ebreak _0282_ _0278_ _1247_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_37_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _1332_ _1341_ _1342_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2885_ _0552_ _0498_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1836_ _1060_ _1277_ _1278_ _1264_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1767_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1698_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _1157_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2319_ _0457_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2249__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3206__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2488__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[2\] net8 net125 u_arbiter.i_wb_cpu_dbus_sel\[0\] net9
+ u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_16_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2117__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2660__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout129_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2670_ _0774_ _0810_ _0813_ _0814_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1621_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3222_ u_cpu.rf_ram_if.wdata0_r\[5\] net39 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input3_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3153_ _0147_ net101 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2104_ u_cpu.cpu.bufreg.lsb\[1\] _0282_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3084_ _0081_ net58 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2035_ u_cpu.rf_ram.i_waddr\[0\] _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout8_I u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2471__B _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2403__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2954__A3 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2868_ _0761_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2799_ _0893_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1819_ _1260_ _1262_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[9\]_SE net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2642__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2881__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2633__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2722_ _0844_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2397__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2653_ _0619_ _0736_ _0597_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2584_ _0609_ _0520_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1604_ u_cpu.rf_ram_if.rtrig0 _1066_ _1072_ _1082_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_47_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout129 net130 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout118 net120 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout107 net109 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3051__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3205_ _0198_ net85 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3136_ _0133_ net119 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3067_ _0064_ net115 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _0225_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _0247_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2624__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2388__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2312__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2615__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2379__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2854__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1814__B1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2305__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2705_ _0835_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2241__S _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2636_ _0779_ _0781_ _0783_ _0455_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2917__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2542__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2567_ _0720_ _0721_ _0612_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2498_ _0537_ _0526_ _0599_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ _0116_ net96 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3097__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2908__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2533__B2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1575__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2524__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2996__S _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2421_ _0587_ _0588_ _0506_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2352_ _0518_ _0521_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2283_ _0430_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[37\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2236__S _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout24_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2212__B1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0227_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1874__I _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2619_ _0543_ _0464_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2373__C _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_scanchain_local.scan_flop\[25\]_SE net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2754__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__B2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[32\]_SI u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3112__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2970_ _0870_ _1009_ _1010_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1921_ _1083_ _1339_ _1352_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1852_ u_cpu.cpu.alu.i_rs1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1783_ u_cpu.rf_ram_if.rdata1\[0\] u_cpu.rf_ram_if.rtrig1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout9 net11 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2404_ _0424_ _0443_ _0572_ _0438_ _0428_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2335_ _0477_ _0505_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2266_ _0432_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2197_ _0385_ _0387_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2520__I1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1711__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2275__I0 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2120_ _0243_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2051_ net2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2953_ u_cpu.cpu.genblk3.csr.mie_mtie _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2966__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1904_ _1331_ u_cpu.rf_ram_if.rdata1\[4\] _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _0616_ _0953_ _0442_ _0594_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ u_cpu.cpu.branch_op _1265_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1766_ _1211_ u_arbiter.o_wb_cpu_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_u_scanchain_local.scan_flop\[0\]_CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3158__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2194__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout91_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ _1154_ _1155_ _1157_ _1158_ u_arbiter.o_wb_cpu_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_103_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2469__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2318_ _0447_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2249_ _1091_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2732__I1 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1999__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2248__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2948__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1620_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_12_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3221_ u_cpu.rf_ram_if.wdata0_r\[4\] net39 u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3152_ _0146_ net99 u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2103_ u_cpu.cpu.bufreg.lsb\[1\] _0282_ _0278_ u_cpu.cpu.bufreg.lsb\[0\] _0312_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3083_ _0080_ net81 u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2034_ _0254_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2308__I _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ _1252_ _0983_ _0986_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1611__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ _0603_ _0611_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2954__A4 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _1084_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0892_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ _1172_ _1197_ _1198_ u_arbiter.o_wb_cpu_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1914__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1678__A1 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2646__C _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1602__A1 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1792__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2837__B _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout141_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2641__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2721_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _0839_
+ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2999__S _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2397__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2652_ _0626_ _0697_ _0568_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2583_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1603_ _1076_ _1080_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout119 net120 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3204_ _0197_ net85 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3135_ _0132_ net108 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3066_ _0063_ net116 u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout54_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2017_ _0225_ _0246_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2482__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ u_arbiter.i_wb_cpu_rdt\[27\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0973_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2388__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2702__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2699__I0 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1823__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1787__I u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[32\] u_arbiter.i_wb_cpu_rdt\[29\] net144 u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ net29 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2000__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__C1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2839__B1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2567__B _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2067__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1814__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1814__B2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2704_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _0833_
+ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ _0502_ _0775_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2321__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2566_ _0689_ _0697_ _0710_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2497_ _0657_ _0469_ _0527_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[6\]_SI u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3118_ _0115_ net76 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3049_ _0046_ net115 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2058__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2908__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2533__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2049__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3041__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout104_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0482_ _0541_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3191__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2351_ _0522_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2282_ _0457_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1997_ _0226_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout17_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2212__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2051__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2618_ _0553_ _0736_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1890__I u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2549_ _0231_ _0677_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2000__B _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2279__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2654__C _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3064__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2136__I _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1920_ u_cpu.rf_ram_if.rdata0\[4\] _1350_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1851_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2745__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1782_ u_cpu.rf_ram.rdata\[0\] _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2403_ _0432_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2334_ _0478_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2265_ _0440_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_113_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2196_ u_arbiter.i_wb_cpu_rdt\[18\] _0386_ _0355_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3087__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2710__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2275__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[21\]_CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1950__A3 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[36\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _0269_ _0255_ _0271_ _1397_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2575__B _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2663__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2415__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2952_ _0997_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2966__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1903_ _1226_ u_cpu.rf_ram.rdata\[4\] _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2883_ _0492_ _0572_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _1045_ _1243_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[20\]_D u_arbiter.i_wb_cpu_rdt\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_1765_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _1210_ _1086_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1696_ u_arbiter.i_wb_cpu_dbus_adr\[15\] _1143_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[15\]_SE net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout84_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2317_ _0425_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2248_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0416_
+ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2179_ _0356_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2654__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_SI u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[11\]_D u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2893__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1696__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2395__B _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2414__I _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[9\]_D u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[62\] u_scanchain_local.module_data_in\[61\] net141 u_arbiter.o_wb_cpu_adr\[24\]
+ net25 u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[38\]_SE net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3220_ u_cpu.rf_ram_if.wdata0_r\[3\] net39 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3151_ _0145_ net101 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2102_ _0281_ _0274_ _0311_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1687__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1931__I0 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2884__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3082_ _0079_ net81 u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2636__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2033_ u_cpu.raddr\[0\] _0248_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3125__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _0983_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1611__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2866_ _0413_ _0521_ _0548_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ _1064_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2260__S _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2797_ _0868_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _1190_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1679_ _1139_ _1140_ _1142_ _1144_ u_arbiter.o_wb_cpu_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1678__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2875__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1850__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1602__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2866__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2837__C _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2618__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3148__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout134_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _0843_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2397__A3 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__I1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2651_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_rdt\[2\] _1094_ _0797_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1602_ u_cpu.cpu.immdec.imm19_12_20\[6\] _1068_ _1069_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_86_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2582_ _0457_ _0547_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3203_ _0196_ net83 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2857__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3134_ _0131_ net108 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3065_ _0062_ net116 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2016_ _0232_ _0245_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2918_ _0974_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2793__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1596__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2849_ _1369_ _1399_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2396__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2699__I1 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2392__C _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1587__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__C2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__B1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2000__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[25\] u_arbiter.i_wb_cpu_rdt\[22\] net131 u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ net16 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_48_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2839__A1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2839__B2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1814__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2703_ _0834_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2634_ _0461_ _0560_ _0766_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ _0523_ _0709_ _0554_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _0523_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3117_ _0114_ net99 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3048_ _0045_ net87 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3007__A1 u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2713__S _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2230__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__C _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2049__A2 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2206__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout91 net93 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout80 net81 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_31_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2221__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2350_ _0523_ _0412_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2281_ _0447_ _0441_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2532__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1996_ u_cpu.cpu.genblk1.align.ctrl_misal _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2212__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _0574_ _0610_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2548_ _0673_ _0701_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2488__B _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2479_ _0590_ _0642_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2279__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2708__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3209__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2451__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3003__I1 u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _1289_ _1291_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1781_ u_cpu.rf_ram.regzero _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2402_ _0528_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2333_ _0491_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2264_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _1090_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2195_ _0342_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2130__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2490__C _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _1084_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3031__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2665__C _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3181__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2735__I0 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2360__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2856__B _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2663__A2 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2147__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2415__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2951_ u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.mstatus_mpie _0980_
+ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ _1332_ _1339_ _1340_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2882_ u_cpu.cpu.immdec.imm11_7\[4\] _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1833_ _1275_ u_cpu.cpu.state.init_done _1057_ _1042_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1764_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1695_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _1142_ _1156_
+ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_63_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__I0 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3054__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2351__A1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout77_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2316_ _0489_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__B _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ _0419_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2178_ _0374_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2721__S _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2717__I0 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2342__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[55\] u_scanchain_local.module_data_in\[54\] net139 u_arbiter.o_wb_cpu_adr\[17\]
+ net24 u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_103_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3077__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2581__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3150_ _0144_ net101 u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3081_ _0078_ net81 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2101_ _1284_ _0286_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2032_ _0253_ _0255_ _0257_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2934_ _1077_ _0984_ _1063_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2865_ _0413_ _0660_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1816_ _1078_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2796_ _0891_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ _1195_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2572__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2340__I _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1678_ u_arbiter.i_wb_cpu_dbus_adr\[11\] _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[20\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[35\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2866__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[0\] net3 net134 u_arbiter.o_wb_cpu_cyc net18 u_cpu.cpu.genblk3.csr.i_mtip
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_114_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2618__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1826__B1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout127_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2650_ _0774_ _0794_ _0795_ _0796_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_12_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ u_cpu.cpu.csr_imm _1067_ _1069_ u_cpu.cpu.immdec.imm24_20\[0\] _1079_ _1080_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_12_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2581_ _0420_ u_arbiter.i_wb_cpu_rdt\[7\] _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2554__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3202_ _0195_ net67 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[12\]_SI u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ _0130_ net108 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3064_ _0061_ net116 u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _1284_ _1057_ _1369_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_24_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1596__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2848_ _0922_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2545__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2779_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0878_ _0880_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2396__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1587__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[35\]_SI u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[18\] u_arbiter.i_wb_cpu_rdt\[15\] net128 u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ net12 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_42_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3115__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2839__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _0833_
+ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2633_ _0489_ _0490_ _0780_ _0686_ _0503_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2564_ _0709_ _0423_ _0561_ _0523_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2495_ _0638_ _0654_ _0655_ _0656_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_29_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3116_ _0113_ net99 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3047_ _0044_ net86 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3007__A2 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2014__B _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2518__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3138__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2206__B1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout81 net85 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout70 net72 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2509__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2280_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _0430_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2748__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1995_ u_cpu.rf_ram_if.rcnt\[0\] _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2616_ _0761_ _0762_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2547_ _0703_ _0594_ _0548_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2488__C _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2478_ u_cpu.cpu.immdec.imm24_20\[2\] _0636_ _0641_ _0486_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1714__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2978__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2433__I _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1780_ _1218_ _1221_ _1222_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2401_ _0477_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _0492_ _0499_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2263_ _0434_ _0435_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2194_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _0375_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1641__A1 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout22_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1978_ _1391_ _1292_ _1393_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1944__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2719__S _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1880__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2253__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2983__I1 u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2360__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1871__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2950_ _0996_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1901_ _1335_ u_cpu.rf_ram_if.rdata1\[3\] _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2881_ _0480_ _0949_ _0950_ _0951_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1832_ u_cpu.cpu.genblk3.csr.o_new_irq _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1763_ _1208_ _1205_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1156_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2315_ _0465_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2351__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2246_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2103__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2177_ u_arbiter.i_wb_cpu_rdt\[12\] _0372_ _0326_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _0373_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[61\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2717__I1 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2878__B1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2342__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2912__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[48\] u_scanchain_local.module_data_in\[47\] net135 u_arbiter.o_wb_cpu_adr\[10\]
+ net19 u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2581__A2 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1771__B _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2100_ _0310_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3080_ _0077_ net79 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2031_ _0256_ u_cpu.rf_ram_if.wen0_r u_cpu.rf_ram_if.rtrig0 _1078_ _0257_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2097__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2933_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2864_ _0600_ _0496_ _0498_ _0537_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1815_ _1060_ _1239_ _1242_ _1245_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2795_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[14\]
+ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1746_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] u_cpu.cpu.ctrl.o_ibus_adr\[25\] u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _1183_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_102_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2021__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ _1101_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2324__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[9\]_SI u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2229_ u_arbiter.i_wb_cpu_rdt\[30\] _0328_ _0400_ u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2088__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2012__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2531__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2866__A3 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1826__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1610__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3044__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1600_ _1052_ _1078_ _1065_ _1067_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2580_ _1092_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2554__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2597__B _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3201_ _0194_ net82 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3132_ _0129_ net108 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3063_ _0060_ net115 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2014_ _1309_ _0242_ _0243_ _1328_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2490__A1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2916_ _0229_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ u_cpu.cpu.immdec.imm11_7\[4\] _0257_ _0259_ u_cpu.rf_ram.i_waddr\[6\] _0922_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2778_ _0881_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1729_ _1177_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3067__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__I _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2472__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2880__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2224__A1 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2701_ _0826_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2171__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2632_ _0549_ _0763_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2563_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _1098_ _0718_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ u_cpu.cpu.immdec.imm24_20\[3\] _0638_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3115_ _0112_ net99 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3046_ _0043_ net114 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[49\]_CLK net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2463__B2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2463__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2014__C _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2518__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2206__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout71 net72 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[30\] u_arbiter.i_wb_cpu_rdt\[27\] net143 u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ net28 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_109_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2445__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1994_ _0224_ _1402_ _1240_ u_arbiter.i_wb_cpu_dbus_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _0549_ _0432_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_u_scanchain_local.scan_flop\[18\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ _0228_ u_arbiter.i_wb_cpu_rdt\[9\] _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_29_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ _0640_ _0636_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3029_ _0011_ net45 u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2436__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1947__B1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2978__A2 u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[32\]_D u_arbiter.i_wb_cpu_rdt\[29\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0492_ _0566_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2589__C _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout102_I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2331_ _0231_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2262_ _0436_ _0437_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_61_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2193_ _0383_ _0384_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2666__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2418__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2969__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3128__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[23\]_D u_arbiter.i_wb_cpu_rdt\[20\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout15_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1977_ _1213_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2529_ _0686_ _0520_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2735__S _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2409__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_D u_arbiter.i_wb_cpu_rdt\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1699__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1900_ _1333_ u_cpu.rf_ram.rdata\[3\] _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ u_cpu.cpu.immdec.imm11_7\[3\] _0923_ _0644_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ u_cpu.cpu.bufreg.lsb\[0\] _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1762_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1693_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1150_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _1155_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2887__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2314_ _0450_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ _0420_ u_arbiter.i_wb_cpu_rdt\[12\] _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2639__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2176_ _0356_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2354__I _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2878__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2878__B2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1608__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2869__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1771__C _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ u_cpu.rf_ram_if.genblk1.wtrig0_r _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2932_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2863_ _0933_ _0935_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2794_ _0890_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1814_ _1056_ _1229_ _1251_ u_cpu.cpu.genblk3.csr.mstatus_mie _1257_ _1258_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1745_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1676_ _1135_ _1125_ _1126_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1780__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__B1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2349__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2228_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2159_ _0356_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1835__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1599__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2812__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__A1 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1826__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2923__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[60\] u_scanchain_local.module_data_in\[59\] net141 u_arbiter.o_wb_cpu_adr\[22\]
+ net25 u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3200_ _0193_ net66 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3131_ _0128_ net108 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2857__A4 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3062_ _0059_ net115 u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2013_ u_arbiter.i_wb_cpu_ack _1101_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2915_ _0972_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2242__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1596__A4 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2846_ _0921_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ _1112_ _0878_ _0880_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1753__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] u_cpu.cpu.ctrl.o_ibus_adr\[22\] _1182_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1659_ _1125_ _1126_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2743__S _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2769__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1867__B _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1744__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3011__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2472__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2224__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3161__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout132_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0832_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1983__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2631_ _0686_ _0611_ _0778_ _0470_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2562_ _0715_ _0716_ _0717_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1735__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2493_ u_cpu.cpu.immdec.imm24_20\[4\] _0474_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2160__A1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3114_ _0111_ net99 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3045_ _0042_ net86 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout45_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2563__S _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2829_ _1195_ _0906_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1726__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3034__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3184__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2206__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1597__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout72 net78 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout50 net52 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1965__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[23\] u_arbiter.i_wb_cpu_rdt\[20\] net131 u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ net16 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2221__B _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2445__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _1039_ _0224_ _1240_ u_arbiter.i_wb_cpu_dbus_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1956__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0598_ _0440_ _0528_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1708__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3057__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _1092_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2476_ u_cpu.cpu.immdec.imm24_20\[1\] _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2133__A1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ _0010_ net40 u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2436__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1947__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2372__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2978__A3 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[33\]_CLK net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[48\]_CLK net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2363__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1705__A4 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _0502_ _0503_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2261_ u_arbiter.i_wb_cpu_rdt\[2\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _0430_
+ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2192_ u_arbiter.i_wb_cpu_rdt\[17\] _0369_ _0370_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2910__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2666__A2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2905__I _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3002__S _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1976_ _1298_ _1279_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2528_ _0418_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2106__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2459_ _0615_ _0622_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_25_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2901__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2657__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2409__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2345__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2648__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[2\]_SE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_19_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1761_ _1139_ _1206_ _1207_ u_arbiter.o_wb_cpu_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2584__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1692_ _1105_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2887__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2313_ _0424_ _0428_ _0442_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_61_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2244_ _0417_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2175_ _0323_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3245__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ _1215_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2327__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2878__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2566__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3118__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2931_ _0980_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2862_ _0689_ _0512_ _0934_ _0486_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2793_ _1145_ _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1813_ _1252_ _1249_ _1253_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2557__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1744_ _1172_ _1193_ _1194_ u_arbiter.o_wb_cpu_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1675_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _1141_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2309__B2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2227_ _0404_ _0406_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _0360_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2365__I _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2089_ _1234_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1599__A2 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2548__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2012__A3 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1619__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2539__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[53\] u_scanchain_local.module_data_in\[52\] net139 u_arbiter.o_wb_cpu_adr\[15\]
+ net23 u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_86_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3130_ _0127_ net106 u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3061_ _0058_ net92 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2012_ _1059_ _1244_ _0241_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2914_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _0967_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2845_ u_cpu.cpu.immdec.imm11_7\[3\] _0257_ _0259_ u_cpu.rf_ram.i_waddr\[5\] _0921_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2776_ _0872_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1727_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _1179_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1658_ _1125_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2163__C1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1589_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_45_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2218__B1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1867__C _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2241__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2941__A1 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ _0687_ _0767_ _0776_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1983__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2561_ _0479_ _0552_ _0712_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2492_ _0484_ _0646_ _0652_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2160__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3113_ _0110_ net100 u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3044_ _0041_ net86 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout38_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2620__B1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2828_ _0910_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2759_ _1213_ _1392_ net2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A3 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout40 net41 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_u_scanchain_local.scan_flop\[41\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout73 net78 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net52 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout62 net68 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout95 net123 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_127_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1965__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[16\] u_arbiter.i_wb_cpu_rdt\[13\] net129 u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ net13 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1632__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1653__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1992_ _1040_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1956__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2613_ _0571_ _0697_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2544_ _0698_ _0700_ _0612_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _0635_ _0638_ _0639_ _0578_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2133__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3027_ _0009_ net42 u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_scanchain_local.scan_flop\[64\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2841__B1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1644__A1 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1947__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2372__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3151__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2484__S _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1635__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2986__I1 u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1938__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1627__I _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2363__A2 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _0430_
+ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2191_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _0375_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1626__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2407__B _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2426__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1975_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1272_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3024__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1929__A2 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3174__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2527_ _0668_ _0683_ _0684_ _0671_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2458_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2389_ _1240_ _0515_ _0559_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1865__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1865__B2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2290__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2345__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[9\] u_arbiter.i_wb_cpu_rdt\[6\] net131 u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ net15 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1856__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3047__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2805__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2281__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1760_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _1143_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2033__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3197__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2584__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ _1153_ u_arbiter.o_wb_cpu_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2312_ _0480_ _0485_ _0487_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2243_ _0226_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3224__D u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2895__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2174_ _0368_ _0371_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2916__I _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1820__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2272__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout20_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1958_ _1106_ _1376_ u_arbiter.o_wb_cpu_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2575__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1889_ _1064_ _1327_ _1330_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2327__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2600__B _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[32\]_CLK net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1838__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[47\]_CLK net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2263__A1 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2566__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2672__S _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _1214_ _1255_ _1249_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2006__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] _0923_ _0934_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2792_ _0889_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1812_ _1213_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1743_ u_arbiter.i_wb_cpu_dbus_adr\[26\] _1190_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3219__D u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2557__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1674_ _1134_ _1136_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2309__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ u_arbiter.i_wb_cpu_rdt\[29\] _0328_ _0405_ u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout68_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2157_ u_arbiter.i_wb_cpu_rdt\[6\] _0324_ _0350_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _0359_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_22_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2088_ _1230_ _0298_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2245__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2381__I _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2181__B1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2539__A2 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[46\] u_scanchain_local.module_data_in\[45\] net135 u_arbiter.o_wb_cpu_adr\[8\]
+ net20 u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3235__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3060_ _0057_ net92 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0238_ _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2913_ _0971_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2415__B _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2844_ _0920_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _0879_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1726_ _1154_ _1178_ _1179_ _1180_ u_arbiter.o_wb_cpu_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1657_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _1113_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1588_ _1037_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2163__B1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ u_arbiter.i_wb_cpu_rdt\[23\] _0386_ _0355_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3189_ _0182_ net86 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2466__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__B2 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2769__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2941__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[2\]_D net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__B1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2457__B2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2457__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2209__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout118_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__B1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ u_cpu.cpu.immdec.imm30_25\[4\] _0706_ _0707_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2491_ _0570_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3112_ _0109_ net100 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3043_ _0040_ net73 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2448__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3232__D u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2620__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2827_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _0906_ _0908_ _1195_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2758_ _0224_ _0863_ _0867_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1709_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _1164_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2689_ _1302_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2439__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A4 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout30 net31 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3080__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout74 net77 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout41 net43 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout52 net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout85 net94 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout96 net98 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__B2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ _1040_ _1402_ _1240_ u_arbiter.i_wb_cpu_dbus_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0703_ _0736_ _0597_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2543_ _0622_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2118__B1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2474_ u_cpu.cpu.immdec.imm24_20\[0\] _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout50_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3026_ _0008_ net42 u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1644__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2841__B2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_scanchain_local.scan_flop\[26\]_D u_arbiter.i_wb_cpu_rdt\[23\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[17\]_D u_arbiter.i_wb_cpu_rdt\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1571__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2190_ _0382_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2426__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1974_ _1390_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1929__A3 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout98_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _0436_ _0499_ _0527_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2457_ _0414_ _0468_ _0519_ _0437_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_u_scanchain_local.scan_flop\[31\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ _0542_ _0552_ _0558_ _0538_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_99_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1865__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3009_ _0019_ net54 u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2290__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2502__B1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2281__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ u_arbiter.i_wb_cpu_dbus_adr\[14\] _1152_ _1087_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout100_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[54\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2311_ _1380_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0415_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2173_ u_arbiter.i_wb_cpu_rdt\[11\] _0369_ _0370_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_0_160 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_fanout13_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3141__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1957_ _1284_ _1370_ _1371_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1888_ _1328_ _1294_ _1329_ _1064_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2509_ _0521_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1838__A2 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2263__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2015__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3014__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3164__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout148_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2860_ _0591_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1811_ u_cpu.cpu.decode.co_ebreak _1049_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2791_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0885_ _0887_ _1145_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1742_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1673_ _1105_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ _0321_ _0316_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2156_ _0325_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2493__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2087_ _1232_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2245__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ u_cpu.rf_ram_if.wdata0_r\[2\] u_cpu.rf_ram_if.wdata1_r\[2\] _1020_ _1021_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2556__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2181__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3037__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[39\] u_scanchain_local.module_data_in\[38\] net132 u_arbiter.o_wb_cpu_adr\[1\]
+ net15 u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _1282_ _0239_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2683__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2912_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _0967_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1600__B _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1986__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2843_ u_cpu.cpu.immdec.imm11_7\[2\] _0257_ _0259_ u_cpu.rf_ram.i_waddr\[4\] _0920_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[31\]_CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2774_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _0878_ _0873_ _1112_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1725_ u_arbiter.i_wb_cpu_dbus_adr\[22\] _1123_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1656_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1587_ _1050_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2163__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2163__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout80_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0357_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3188_ _0181_ net59 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2139_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _0320_ _0316_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2218__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1977__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__B2 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1901__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2209__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1968__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3202__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ _0575_ _0648_ _0650_ _0651_ _0483_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2393__B2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3111_ _0108_ net73 u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3042_ _0039_ net75 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2826_ _0909_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2620__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2757_ _0863_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2688_ _0825_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1708_ _1154_ _1164_ _1165_ _1166_ u_arbiter.o_wb_cpu_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1639_ _1106_ _1110_ _1111_ u_arbiter.o_wb_cpu_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2439__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout20 net21 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3225__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout42 net43 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout53 net62 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout86 net88 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout75 net77 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout97 net98 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_13_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2375__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2297__I _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1990_ u_cpu.cpu.bne_or_bge _1039_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2989__I0 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout130_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2760__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2611_ _0759_ _0752_ _0760_ _0564_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2542_ _0600_ _0613_ _0614_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2366__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[18\]_SI u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2118__B2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2118__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2473_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2669__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3248__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ _0007_ net48 u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2841__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout43_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2809_ _0868_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2357__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2109__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[21\] u_arbiter.i_wb_cpu_rdt\[18\] net130 u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ net12 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_26_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1973_ _1378_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2587__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2339__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2525_ _0482_ _0626_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2456_ _0611_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2511__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _0517_ _0557_ _0491_ _0552_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3008_ _0259_ _1032_ _1033_ _1034_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_25_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2578__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2750__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2502__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1856__A3 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2805__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[69\] u_scanchain_local.module_data_in\[68\] net147 u_arbiter.o_wb_cpu_adr\[31\]
+ net30 u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_15_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3093__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1654__I _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2310_ _0478_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2241_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _0417_
+ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0325_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1829__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2434__B _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _1373_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2280__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1765__S _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1887_ _1274_ _1285_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1783__A2 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2508_ _0542_ _0613_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2439_ _0570_ _0455_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2015__A3 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2971__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1810_ u_cpu.cpu.decode.op21 _1044_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_SE net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2790_ _0888_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1741_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _1185_ _1183_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1672_ _1133_ _1138_ u_arbiter.o_wb_cpu_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2962__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3411_ u_scanchain_local.data_out net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2224_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _0400_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2155_ _0354_ _0358_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2086_ _1242_ _1277_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ u_cpu.rf_ram_if.genblk1.wtrig0_r _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1939_ u_cpu.rf_ram.i_waddr\[3\] _1362_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1756__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2556__I1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2181__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2157__C1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1932__I _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2763__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _0970_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1600__C _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[7] u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1986__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2842_ _0919_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2773_ _0869_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2235__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ _1176_ _1177_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1655_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1586_ _1056_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2163__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout73_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2207_ _0393_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3187_ _0180_ net51 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2138_ _0320_ _0235_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[67\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2710__I1 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2069_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1977__A2 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3154__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1665__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2583__I _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1968__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[51\] u_scanchain_local.module_data_in\[50\] net136 u_arbiter.o_wb_cpu_adr\[13\]
+ net19 u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2378__C1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.out_flop u_scanchain_local.module_data_in\[69\] net31 u_scanchain_local.data_out_i
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_64_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3110_ _0107_ net70 u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3041_ _0038_ net72 u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2081__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _0906_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2756_ _0858_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3177__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2384__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2687_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _1378_ _0825_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1707_ u_arbiter.i_wb_cpu_dbus_adr\[18\] _1123_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1638_ u_arbiter.i_wb_cpu_dbus_adr\[4\] _1103_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1569_ _1046_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1572__I u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1895__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3239_ u_cpu.cpu.o_wen0 net56 u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2695__I0 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout10 net11 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout21 net26 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout32 net33 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout54 net61 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout43 net44 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout65 net67 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net102 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout76 net78 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2375__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[30\]_CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2835__B1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2989__I1 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ u_cpu.cpu.csr_imm _0644_ _0755_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2541_ _0413_ _0697_ _0541_ _0609_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2366__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2472_ _0570_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2118__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1877__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1629__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ _0027_ net56 u_cpu.rf_ram.i_waddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout36_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2054__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2808_ _0898_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2357__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2739_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _0851_
+ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2293__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2348__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1571__A3 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[14\] u_arbiter.i_wb_cpu_rdt\[11\] net128 u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ net12 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_26_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2284__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2036__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1972_ _1379_ _1383_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2587__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2524_ _0634_ _0682_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2455_ _0616_ _0617_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2386_ _0481_ _0464_ _0553_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2511__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ u_cpu.rf_ram.i_wdata\[7\] _0263_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2502__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2266__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2240_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2171_ _0342_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_D[7] u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2009__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ _1264_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1886_ _1042_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2980__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ _0664_ _0667_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2438_ _0594_ _0602_ _0603_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1580__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2369_ _0519_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2971__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2184__B1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[7\] u_arbiter.i_wb_cpu_rdt\[4\] net132 u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ net15 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_130_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1740_ _1172_ _1189_ _1191_ u_arbiter.o_wb_cpu_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2411__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ _1134_ _1136_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3410_ u_scanchain_local.clk_out net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2223_ _0403_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2154_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0355_ _0357_ _0241_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2085_ _1317_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ _1019_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1938_ _1080_ _1361_ _1363_ u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1869_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2166__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3083__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2157__B1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2157__C2 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[5\]_D u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1683__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2880__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2910_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _0967_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2632__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_A[6] u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2841_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _0869_ _0872_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2772_ _0877_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1723_ _1176_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2148__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ _1101_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1585_ _1057_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2206_ u_arbiter.i_wb_cpu_rdt\[22\] _0372_ _0359_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _0373_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_41_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3186_ _0179_ net57 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2137_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2871__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2068_ _0272_ _0273_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2623__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[11\]_SE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2862__B2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2862__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2614__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2378__C2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[44\] u_scanchain_local.module_data_in\[43\] net138 u_arbiter.o_wb_cpu_adr\[6\]
+ net22 u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__S _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3040_ _0037_ net74 u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2853__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2853__B2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__B2 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2081__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2824_ _0871_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2755_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _1400_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2686_ _0824_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1706_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _1160_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _1165_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1637_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1568_ u_cpu.cpu.bne_or_bge _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2541__B1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3238_ u_cpu.cpu.o_wdata1 net55 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3169_ _0163_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[29\]_D u_arbiter.i_wb_cpu_rdt\[26\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2695__I1 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout11 net14 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout22 net26 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout33 net34 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2072__A2 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout55 net61 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout44 net69 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_52_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout88 net93 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout77 net78 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout99 net100 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout66 net67 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3121__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1583__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1638__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2540_ _0468_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2771__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1673__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[57\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1574__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ _0297_ _1377_ _1044_ _1214_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_64_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2523__B1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1629__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3023_ _0026_ net56 u_cpu.rf_ram.i_waddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__C _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout29_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3144__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _0892_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2738_ _0853_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1565__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ u_cpu.cpu.immdec.imm19_12_20\[8\] _0751_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2514__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2293__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2045__A2 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3017__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2284__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ _1384_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1795__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2499__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ u_cpu.cpu.immdec.imm30_25\[1\] _0678_ _0679_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2454_ _0411_ _0619_ _0598_ _0522_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2385_ _0412_ _0537_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3006_ _0256_ u_cpu.rf_ram_if.wdata1_r\[7\] _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[59\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2112__I _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1951__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _0361_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1701__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__S _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2257__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_D[6] u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2009__A2 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1954_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1885_ _1267_ _1294_ _1310_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout96_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ u_cpu.cpu.immdec.imm24_20\[4\] _0637_ _0661_ _0512_ _0666_ _0667_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_44_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ _0436_ _0571_ _0502_ _0593_ _0575_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ _0471_ _0469_ _0483_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2299_ _0475_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2971__A3 u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2184__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3205__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2107__I _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2411__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1670_ _1134_ _1136_ _1105_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ u_arbiter.i_wb_cpu_rdt\[28\] _0342_ _0359_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _0356_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2478__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2153_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2084_ u_cpu.cpu.ctrl.i_jump _0286_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1989__A1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout11_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2986_ _1018_ u_cpu.rf_ram.i_wdata\[1\] _0263_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1937_ u_cpu.rf_ram.i_waddr\[2\] _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1868_ u_cpu.cpu.state.o_cnt_r\[1\] _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2166__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ u_cpu.cpu.decode.co_mem_word _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2469__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2713__I0 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3228__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2157__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[8\]_SE net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout146_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[5] u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2840_ _0916_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2771_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0870_ _0873_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1722_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] u_cpu.cpu.ctrl.o_ibus_adr\[20\] u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _1164_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_8_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1653_ _1106_ _1121_ _1122_ u_arbiter.o_wb_cpu_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2148__B2 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2148__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1584_ _1058_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2205_ _0391_ _0392_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2320__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ _0178_ net64 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2136_ _0323_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout59_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2871__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2067_ _0281_ _0284_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2969_ u_cpu.cpu.state.ibus_cyc _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2387__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2139__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3050__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2311__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2862__A2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2614__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2378__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__B2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[37\] u_scanchain_local.module_data_in\[36\] net145 u_arbiter.i_wb_cpu_dbus_dat\[31\]
+ net27 u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__I _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2550__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2853__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2991__S _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2081__A3 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2823_ _0907_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2754_ _1274_ _0863_ _0864_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1705_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _1157_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _1378_ _0824_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1636_ _1098_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _1096_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1592__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3073__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1567_ u_cpu.cpu.decode.co_mem_word _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2541__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2541__B2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2030__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3237_ u_cpu.rf_ram_if.wdata1_r\[7\] net45 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3168_ _0162_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2119_ _0319_ _0322_ _0327_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3099_ _0096_ net57 u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout12 net13 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout34 u_scanchain_local.clk net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout23 net25 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout45 net53 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout56 net60 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout89 net91 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout78 net95 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout67 net68 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2835__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2115__I _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2220__B1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1954__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ u_cpu.cpu.immdec.imm24_20\[1\] _0479_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2986__S _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2785__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3022_ _0025_ net46 u_cpu.rf_ram.i_waddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2806_ _0897_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2737_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _0851_
+ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2762__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2668_ _1373_ _0727_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1619_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_47_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2599_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2514__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2628__C _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2753__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2554__B _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1949__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _1309_ _1225_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[24\]_SE net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ _0675_ _0681_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2453_ _0420_ u_arbiter.i_wb_cpu_rdt\[10\] _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2384_ _0523_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2448__C _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3005_ _0265_ u_cpu.cpu.o_wdata0 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout41_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1786__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1769__I _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_D[5] u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserv_0_153 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ _1263_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2965__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1884_ _1316_ _1318_ _1258_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2505_ _0637_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2436_ _0435_ _0541_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1940__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout89_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2367_ _0444_ _0507_ _0512_ _0537_ _0539_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2298_ _0297_ _0473_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1589__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1759__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2956__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2184__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[67\] u_scanchain_local.module_data_in\[66\] net147 u_arbiter.o_wb_cpu_adr\[29\]
+ net30 u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2947__A1 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _0399_ _0400_ _0402_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2994__S _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0349_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2083_ _0293_ _0295_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[43\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__S _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2985_ u_cpu.rf_ram_if.wdata0_r\[1\] u_cpu.rf_ram_if.wdata1_r\[1\] _0265_ _1018_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2938__B2 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2938__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1936_ _1357_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_15_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1867_ _1297_ _1308_ _1309_ _1278_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1798_ _1240_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2166__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _0503_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2636__C _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2929__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__B2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1601__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2157__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1840__A1 u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_A[4] u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ _0876_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout139_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2989__S _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ u_arbiter.i_wb_cpu_dbus_adr\[7\] _1115_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2148__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2788__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1583_ u_cpu.cpu.decode.op21 _1053_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_119_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2204_ u_arbiter.i_wb_cpu_rdt\[21\] _0386_ _0355_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3184_ _0177_ net66 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2135_ u_arbiter.i_wb_cpu_rdt\[3\] _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2320__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2066_ _0282_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2968_ _0653_ _0285_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1919_ _1083_ _1337_ _1351_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2899_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _0961_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1898__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2847__B1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2311__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2075__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2401__I _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2550__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2557__B _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2861__I0 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2822_ _1185_ _0906_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2753_ _1040_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _1124_ _1162_ _1163_ u_arbiter.o_wb_cpu_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2684_ _0823_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1635_ _1106_ _1107_ _1108_ u_arbiter.o_wb_cpu_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1566_ u_cpu.cpu.csr_d_sel _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2541__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout71_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3236_ u_cpu.rf_ram_if.wdata1_r\[6\] net40 u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3167_ _0161_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2118_ u_arbiter.i_wb_cpu_rdt\[0\] _0324_ _0326_ _1321_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3098_ _0095_ net66 u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2057__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ _0256_ u_cpu.cpu.immdec.imm11_7\[1\] _0254_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_78_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout13 net14 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout35 u_arbiter.i_wb_cpu_dbus_dat\[1\] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout24 net25 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout46 net53 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout68 net69 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout57 net60 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout79 net81 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1583__A3 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2048__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2220__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2771__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3021_ _0024_ net46 u_cpu.rf_ram.i_waddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2306__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2805_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _0892_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3040__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2736_ _0852_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2211__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2667_ _0532_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1618_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_47_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3190__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2598_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2514__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3219_ u_cpu.rf_ram_if.wdata0_r\[2\] net37 u_cpu.rf_ram_if.wdata0_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2450__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3063__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2441__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2997__S _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ u_cpu.cpu.immdec.imm30_25\[0\] _0678_ _0679_ u_cpu.cpu.immdec.imm30_25\[1\]
+ _0580_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_100_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1952__B1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2452_ _0417_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2383_ _0522_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 io_in[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3004_ _1031_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2745__B _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2680__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2237__S _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2432__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _0839_
+ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3086__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2671__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__B1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1785__I0 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[12\] u_arbiter.i_wb_cpu_rdt\[9\] net125 u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ net9 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_D[4] u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__B _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserv_0_154 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ _1244_ _1040_ _1048_ _1039_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1883_ _0037_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2520__S _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2504_ u_cpu.cpu.immdec.imm30_25\[0\] _0532_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2435_ _0596_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2366_ _1373_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2297_ _0231_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2653__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[10\]_D u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2892__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_D u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3101__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2220_ u_arbiter.i_wb_cpu_rdt\[27\] _0324_ _0350_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2151_ _0325_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2883__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2082_ _0028_ _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__B _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__A1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2984_ _1017_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2938__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1935_ _1357_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__2314__I _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ _1043_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1797_ _1047_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_u_scanchain_local.scan_flop\[37\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2418_ _0582_ _0584_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2349_ _0411_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2874__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2874__B2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3124__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2929__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__A2 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2894__I _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[5\] u_arbiter.i_wb_cpu_rdt\[2\] net126 u_arbiter.i_wb_cpu_dbus_sel\[3\]
+ net10 u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2865__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2093__A2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_A[3] u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ _1172_ _1174_ _1175_ u_arbiter.o_wb_cpu_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _1118_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1582_ _1059_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2203_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _0357_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3183_ _0176_ net57 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2856__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2134_ _0340_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2065_ _0278_ _0277_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2608__B2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3147__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2084__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2967_ _0272_ u_cpu.cpu.genblk3.csr.timer_irq_r _0820_ _1008_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_13_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _0963_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1595__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ u_cpu.rf_ram_if.rdata0\[3\] _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1849_ _1273_ _1288_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2847__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2647__C _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2663__B _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1793__I u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[42\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2557__C _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[57\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1813__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2861__I1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2821_ _0868_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ _1285_ _0233_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2774__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1703_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _1147_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2683_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _1378_ _0823_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ u_arbiter.i_wb_cpu_dbus_adr\[3\] _1103_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1565_ _1042_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3235_ u_cpu.rf_ram_if.wdata1_r\[5\] net40 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ _0160_ net104 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2117_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2039__I _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3097_ _0094_ net66 u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2048_ _0256_ _1051_ _1268_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_93_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1878__I u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout14 net17 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout25 net26 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout36 net38 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout47 net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout69 net124 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3006__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout58 net60 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2765__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1740__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2220__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[42\] u_scanchain_local.module_data_in\[41\] net137 u_arbiter.o_wb_cpu_adr\[4\]
+ net21 u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1731__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3020_ _0023_ net50 u_cpu.rf_ram.i_waddr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1798__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2804_ _0896_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2211__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2735_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _0851_
+ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2666_ _1328_ u_cpu.cpu.immdec.imm24_20\[0\] _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1970__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ _1214_ _0749_ _0230_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3218_ u_cpu.rf_ram_if.wdata0_r\[1\] net36 u_cpu.rf_ram_if.wdata0_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3149_ _0143_ net101 u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2450__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3002__I1 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3208__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2441__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2520_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_rdt\[9\] _1095_ _0680_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1952__B2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2451_ _0422_ _0493_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1704__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2382_ _0422_ _0495_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput4 io_in[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3003_ _1030_ u_cpu.rf_ram.i_wdata\[6\] _1022_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2317__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout27_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2196__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2718_ _0842_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2052__I _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ u_cpu.cpu.immdec.imm19_12_20\[6\] _0751_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1785__I1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[3] u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3030__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2662__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserv_0_155 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2137__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3180__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1882_ _1236_ _1323_ _1317_ _1264_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2503_ _0606_ _0659_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2434_ _0597_ _0599_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ _0230_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2296_ _0424_ _0444_ _0456_ _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2475__C _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2653__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2047__I u_cpu.rf_ram.i_waddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1886__I _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3053__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2580__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2332__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ u_arbiter.i_wb_cpu_rdt\[5\] _0343_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2081_ _1373_ _1374_ _1371_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2635__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ _1016_ u_cpu.rf_ram.i_wdata\[0\] _0263_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1934_ _1360_ u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2399__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1865_ _1039_ _1302_ _1305_ _1236_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1796_ _1046_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3076__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2571__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2417_ _0527_ _0481_ _0572_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2348_ _0448_ _0457_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2874__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2279_ _0445_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2706__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2865__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_A[2] u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1840__A3 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3099__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1650_ _1117_ _1119_ _1120_ u_arbiter.o_wb_cpu_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1581_ u_cpu.cpu.decode.co_mem_word u_cpu.cpu.bne_or_bge _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2202_ _0390_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3182_ _0013_ net79 u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2133_ u_arbiter.i_wb_cpu_rdt\[2\] _0328_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ u_cpu.cpu.mem_bytecnt\[1\] _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2966_ _1058_ _0286_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2897_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _0961_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1917_ _1067_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2261__S _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1848_ _1290_ _1249_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1595__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2919__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2060__I _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1779_ u_cpu.cpu.bufreg2.i_cnt_done u_cpu.cpu.immdec.imm31 _1223_ _1224_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[11\]_SI u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2838__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[27\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout144_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _0905_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2751_ u_cpu.cpu.state.o_cnt_r\[1\] _1290_ _1249_ _0233_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1984__I _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2682_ _0822_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1702_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _1160_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1633_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _1099_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2526__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1564_ u_cpu.cpu.decode.opcode\[2\] _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3114__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3234_ u_cpu.rf_ram_if.wdata1_r\[4\] net39 u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3165_ _0159_ net104 u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2116_ _0323_ _0315_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout57_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3096_ _0093_ net80 u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2047_ u_cpu.rf_ram.i_waddr\[3\] _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout15 net17 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout26 net33 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__B1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout37 net38 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3006__A2 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout48 net52 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout59 net60 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_104_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2214__C2 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2214__B1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _0994_ u_cpu.cpu.genblk3.csr.mcause31 _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2765__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2765__B2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2517__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1879__I0 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2048__A3 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2508__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[35\] u_scanchain_local.module_data_in\[34\] net145 u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ net27 u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1798__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2803_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _0892_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2747__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2603__I _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ _1302_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2665_ _0657_ _0764_ _0806_ _0471_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_47_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2759__B net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1970__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1616_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ _1223_ _1266_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2478__C _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3217_ _0209_ net114 u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3148_ _0142_ net114 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3079_ _0076_ net59 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[41\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[56\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2388__C _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2977__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout107_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1952__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ _0496_ _0494_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2381_ _0505_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3002_ u_cpu.rf_ram_if.wdata0_r\[6\] u_cpu.rf_ram_if.wdata1_r\[6\] _1020_ _1030_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2968__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2196__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2717_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _0839_
+ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2991__I1 u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2648_ u_cpu.cpu.immdec.imm19_12_20\[7\] _0514_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2579_ _0582_ _0731_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2743__I1 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2259__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2959__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2187__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2431__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_D[2] u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xserv_0_156 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ u_cpu.cpu.state.o_cnt_r\[1\] _1290_ _1246_ u_cpu.cpu.state.o_cnt_r\[2\] _1369_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1881_ _1243_ _1319_ _1320_ _1323_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1622__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2153__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__I _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2502_ _0582_ _0537_ _0587_ _0662_ _0504_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ _0435_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2364_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ _0464_ _0469_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2810__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2063__I _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2413__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1916__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[60\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2801__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1604__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2701__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2080_ _1077_ _0286_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2096__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__I _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2592__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2982_ u_cpu.rf_ram_if.wdata0_r\[0\] u_cpu.rf_ram_if.wdata1_r\[0\] _0265_ _1016_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ u_cpu.raddr\[1\] u_cpu.rf_ram.i_waddr\[1\] _1358_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2399__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1864_ _1059_ _1244_ u_cpu.cpu.alu.cmp_r _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_102_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1795_ _1236_ _1232_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2020__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2571__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2416_ _0481_ _0583_ _0567_ _0489_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout87_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2347_ _0468_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2278_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2087__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1834__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3020__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[1] u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[65\] u_scanchain_local.module_data_in\[64\] net147 u_arbiter.o_wb_cpu_adr\[27\]
+ net30 u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2250__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _1045_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2002__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3250_ _0223_ net46 u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2201_ u_arbiter.i_wb_cpu_rdt\[20\] _0372_ _0359_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _0373_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_117_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3181_ _0175_ net50 u_cpu.rf_ram.i_waddr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2132_ _0335_ _0337_ _0321_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0272_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1816__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2965_ _0673_ _1007_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2896_ _0962_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1916_ _1083_ _1334_ _1349_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1847_ u_cpu.cpu.state.o_cnt_r\[0\] _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_15_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3193__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1778_ u_cpu.cpu.branch_op u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.csr_d_sel _1223_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2497__B _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2717__S _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1807__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2627__S _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2854__C _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3066__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2471__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2750_ _1285_ _0858_ _0861_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout137_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2681_ u_arbiter.i_wb_cpu_dbus_adr\[2\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _1378_ _0822_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1701_ _1154_ _1159_ _1160_ _1161_ u_arbiter.o_wb_cpu_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1563_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3233_ u_cpu.rf_ram_if.wdata1_r\[3\] net37 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3164_ _0158_ net103 u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2115_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3095_ _0092_ net80 u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2046_ _0255_ _0267_ _0268_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout16 net17 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout27 net29 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2462__B2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout38 net43 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout49 net52 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2214__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2948_ _0273_ _1255_ _1261_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2765__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2879_ u_cpu.cpu.immdec.imm11_7\[4\] _1370_ _1399_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1879__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2910__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[28\] u_arbiter.i_wb_cpu_rdt\[25\] net143 u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ net28 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_7_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2156__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2444__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2802_ _0895_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2733_ _0850_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2747__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2664_ _0538_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1970__A3 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1615_ u_cpu.cpu.genblk1.align.ctrl_misal _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2595_ _1309_ _1380_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3216_ _0017_ net48 u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3147_ _0141_ net100 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ _0075_ net66 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2029_ _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[17\]_SE net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[31\]_D u_arbiter.i_wb_cpu_rdt\[28\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2380_ _1241_ _0515_ _0551_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3001_ _1029_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2665__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2665__B2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__A1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2968__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[22\]_D u_arbiter.i_wb_cpu_rdt\[19\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_2716_ _0841_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2647_ _0484_ _0788_ _0790_ _0793_ _0653_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2578_ _0627_ _0442_ _0497_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2656__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2259__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2408__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3127__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2959__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[13\]_D u_arbiter.i_wb_cpu_rdt\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1698__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[1] u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2647__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1870__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xserv_0_157 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _1243_ _1320_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2501_ _0657_ _0529_ _0660_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2432_ _0598_ _0463_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2363_ _0228_ u_arbiter.i_wb_cpu_rdt\[6\] _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2886__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[40\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2294_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2638__A1 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout32_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2280__S _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2413__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2877__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A1 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1604__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[10\] u_arbiter.i_wb_cpu_rdt\[7\] net128 u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ net12 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_79_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2981_ _0281_ _0232_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1932_ _1359_ u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1863_ _1290_ _1248_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1794_ _1236_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2113__B _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2415_ _0496_ _0494_ _0465_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2859__B2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2346_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2277_ _0448_ _0451_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1834__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2795__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_A[0] u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2250__A2 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2712__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[58\] u_scanchain_local.module_data_in\[57\] net140 u_arbiter.o_wb_cpu_adr\[20\]
+ net24 u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2002__A2 u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1761__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2200_ _0388_ _0389_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3180_ _0174_ net50 u_cpu.rf_ram.i_waddr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2159__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2131_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _0331_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2062_ _0278_ _0277_ _0280_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1998__I _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1816__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2964_ u_cpu.cpu.ctrl.i_iscomp _0480_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1915_ u_cpu.rf_ram_if.rdata0\[2\] _1347_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _1273_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1777_ u_arbiter.i_wb_cpu_dbus_we _1220_ u_cpu.cpu.immdec.imm24_20\[0\] _1222_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2069__I _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ _0453_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_61_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1807__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2465__C1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2232__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1743__A1 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2908__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[3\] u_arbiter.i_wb_cpu_rdt\[0\] net125 u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ net9 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2471__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1700_ u_arbiter.i_wb_cpu_dbus_adr\[16\] _1143_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ _1396_ _0307_ _0821_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1631_ _1102_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1562_ u_cpu.cpu.branch_op _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3232_ u_cpu.rf_ram_if.wdata1_r\[2\] net36 u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input4_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ _0157_ net103 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2114_ net8 _1101_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3094_ _0091_ net79 u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3010__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ u_cpu.rf_ram.i_waddr\[2\] _0263_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout28 net29 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout17 net18 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2462__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3160__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout39 net41 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2214__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout9_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2947_ _1275_ _1260_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1973__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2878_ _0529_ _0587_ _0554_ _0471_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1725__A1 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2150__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1879__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A2 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2141__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3033__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3183__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2444__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2801_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _0892_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2172__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2732_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _0845_
+ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _1098_ u_arbiter.i_wb_cpu_rdt\[19\] _0483_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1614_ _1089_ u_arbiter.o_wb_cpu_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1707__A1 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2594_ _0745_ _0746_ _0747_ _1396_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2380__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3215_ _0208_ net71 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3146_ _0015_ net75 u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout62_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3077_ _0074_ net58 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2028_ u_cpu.rf_ram_if.genblk1.wtrig0_r u_cpu.rf_ram_if.wen1_r _1038_ u_cpu.rf_ram_if.wen0_r
+ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2199__A1 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3056__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2674__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2921__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[40\] u_scanchain_local.module_data_in\[39\] net145 u_arbiter.o_wb_cpu_adr\[2\]
+ net27 u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2362__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2114__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3000_ _1028_ u_cpu.rf_ram.i_wdata\[5\] _1022_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2417__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2715_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _0839_
+ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2646_ _0703_ _0765_ _0792_ _0594_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2577_ _0419_ _0609_ _0443_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2105__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2656__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3129_ _0126_ net106 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2741__S _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2592__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2719__I0 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_D[0] u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2647__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xserv_0_158 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout112_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2500_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _0592_ _0661_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2431_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0417_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2335__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2362_ _1092_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2886__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2293_ _0450_ _0452_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2638__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1861__A3 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[1\]_SE net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout25_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2574__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2326__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2629_ _0686_ _0522_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[14\]_SI u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__A2 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2980_ _1356_ _1362_ _0255_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1931_ u_cpu.raddr\[0\] u_cpu.rf_ram.i_waddr\[0\] _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ u_cpu.cpu.bne_or_bge _1303_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1793_ u_cpu.cpu.csr_imm _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3117__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2414_ _0452_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2345_ _0493_ _0501_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2276_ _0425_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2795__B2 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[54\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2130_ _0316_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[69\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2061_ _0278_ _0277_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2175__I _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2226__B1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2963_ _1003_ _1004_ _1005_ _1006_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_128_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _1083_ _1227_ _1348_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2894_ _0229_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3000__S _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1845_ _1274_ _1285_ _1267_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_15_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2529__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1776_ u_arbiter.i_wb_cpu_dbus_we _1219_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_102_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1752__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2328_ _0425_ _0452_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2259_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] _1090_
+ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1807__A3 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__C2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__B1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2085__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1743__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2723__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2759__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _1097_ _1100_ _1104_ u_arbiter.o_wb_cpu_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1561_ _1039_ _1040_ u_arbiter.i_wb_cpu_dbus_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1734__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3231_ u_cpu.rf_ram_if.wdata1_r\[1\] net36 u_cpu.rf_ram_if.wdata1_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3162_ _0156_ net103 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2113_ net35 _0320_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3093_ _0090_ net79 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2044_ _0265_ u_cpu.cpu.immdec.imm11_7\[0\] _1261_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2298__I0 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout29 net32 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout18 net34 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2946_ _0992_ _0983_ _0993_ _1260_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2877_ _0709_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1828_ _1220_ _1269_ _1270_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1693__B u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1725__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2150__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1879__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__A1 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1964__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2919__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2141__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1652__A1 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout142_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2800_ _0871_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[40\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0849_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2662_ _1094_ _0341_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xu_scanchain_local.output_buffers\[2\] u_scanchain_local.data_out_i u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1613_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _1086_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2593_ u_cpu.cpu.immdec.imm7 _0591_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1707__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2380__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3214_ _0207_ net59 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3145_ _0016_ net75 u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout55_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3076_ _0073_ net58 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2027_ u_cpu.rf_ram.i_waddr\[7\] _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2691__I0 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2199__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2929_ _1218_ _1064_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2994__I1 u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1946__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2739__S _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1882__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_SE net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1937__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1617__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[33\] u_arbiter.i_wb_cpu_rdt\[30\] net144 u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ net29 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_68_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2362__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2876__C _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3150__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2114__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0840_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2050__B2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2132__B _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2645_ _0761_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2576_ _0723_ _0724_ _0730_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1864__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3128_ _0125_ net105 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3059_ _0056_ net91 u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2821__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3023__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2592__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3173__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2268__I _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1855__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xserv_0_159 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout105_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _0516_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2887__B _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2335__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ _1377_ _0515_ _0534_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2292_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2099__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3003__S _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3046__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout18_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3196__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2023__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2326__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _0436_ _0613_ _0458_ _0542_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2559_ _0673_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1837__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2037__B u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2262__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2927__S _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3069__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1930_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1861_ _1243_ _1232_ _1230_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2461__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1792_ _1045_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1805__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2410__B _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2413_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _1098_ _0581_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2344_ _0459_ _0462_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2275_ u_arbiter.i_wb_cpu_rdt\[1\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _0416_
+ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2492__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2244__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__I _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2547__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3211__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__B2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2538__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2884__C _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _1085_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2474__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2226__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2962_ u_cpu.cpu.genblk3.csr.mstatus_mie _1003_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1913_ u_cpu.rf_ram_if.rdata0\[1\] _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2893_ _0281_ _0960_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1844_ u_cpu.cpu.mem_bytecnt\[1\] _1286_ _1267_ _1225_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_15_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2529__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1775_ u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.decode.opcode\[0\] u_cpu.cpu.decode.opcode\[1\]
+ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2140__B _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout85_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2327_ _0465_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2258_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _0416_
+ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2189_ u_arbiter.i_wb_cpu_rdt\[16\] _0372_ _0326_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _0373_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__1807__A4 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__B2 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2217__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[1\]_D u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2456__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2208__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2759__A2 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[63\] u_scanchain_local.module_data_in\[62\] net142 u_arbiter.o_wb_cpu_adr\[25\]
+ net25 u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1560_ u_cpu.cpu.bufreg.lsb\[1\] _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2392__B1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3230_ _0213_ net48 u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3161_ _0155_ net102 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2112_ _0243_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3092_ _0089_ net64 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3222__D u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ _1052_ _1261_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout19 net21 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2945_ _1268_ _1062_ _0982_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2876_ _0582_ _0697_ _0944_ _0575_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1827_ _1265_ u_cpu.cpu.decode.opcode\[1\] _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1758_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _1196_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1689_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1150_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2438__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2824__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1661__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[53\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[68\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1884__B _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2374__B1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2429__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2734__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[34\]_D u_arbiter.i_wb_cpu_rdt\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _0845_
+ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout135_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__B2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2601__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2661_ _0568_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1612_ _1088_ u_arbiter.o_wb_cpu_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2592_ _1370_ _0727_ _0644_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3213_ _0206_ net70 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2668__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3144_ _0140_ net86 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3075_ _0072_ net113 u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2026_ _0246_ _0252_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1969__B _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout48_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2691__I1 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[25\]_D u_arbiter.i_wb_cpu_rdt\[22\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0979_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2859_ _0929_ _0930_ _0931_ _0587_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1634__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[16\]_D u_arbiter.i_wb_cpu_rdt\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[26\] u_arbiter.i_wb_cpu_rdt\[23\] net143 u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ net28 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1570__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2713_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _0839_
+ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2050__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2644_ _0599_ _0767_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2889__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2575_ u_cpu.cpu.immdec.imm7 _1382_ _0679_ _0729_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2338__B1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1561__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3127_ _0124_ net105 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3058_ _0055_ net89 u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2009_ _1218_ _1392_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[30\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__B1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2032__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0517_ _0526_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2291_ _0465_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A2 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A1 u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2627_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _1093_ _0775_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[53\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2558_ _0612_ _0711_ _0713_ _0490_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2489_ _0543_ _0610_ _0574_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2798__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3140__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1860_ _1295_ _1230_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2005__A2 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1791_ _1214_ _1216_ _1235_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2412_ _0510_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2343_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2274_ _0450_ _0427_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3013__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2492__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout30_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__A3 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1989_ _1397_ _1401_ _1396_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1887__B _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1994__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2511__B _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3036__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2226__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ u_cpu.cpu.genblk3.csr.mstatus_mpie _1050_ _1397_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1912_ _1068_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2892_ _1095_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1985__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1774_ u_cpu.cpu.immdec.imm11_7\[0\] _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2326_ _0227_ u_arbiter.i_wb_cpu_rdt\[15\] _0500_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_fanout78_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2257_ _0417_ _0341_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2188_ _0380_ _0381_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2465__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2217__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3059__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1900__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2208__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[56\] u_scanchain_local.module_data_in\[55\] net139 u_arbiter.o_wb_cpu_adr\[18\]
+ net23 u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2392__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2144__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3160_ _0154_ net96 u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2111_ _0234_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3091_ _0088_ net47 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2042_ u_cpu.rf_ram_if.genblk1.wtrig0_r _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__B _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1958__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2944_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2875_ _0925_ _0942_ _0946_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3201__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _1041_ _1215_ _1268_ _1053_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1757_ _1139_ _1203_ _1204_ u_arbiter.o_wb_cpu_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1688_ _1139_ _1149_ _1150_ _1151_ u_arbiter.o_wb_cpu_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ _0482_ _0484_ _0469_ _0471_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A2 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1884__C _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2061__B _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2374__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2374__B2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2126__A1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2677__A2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2921__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[1\] u_cpu.cpu.genblk3.csr.i_mtip net134 u_arbiter.o_wb_cpu_we
+ net18 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0657_ _0737_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1611_ _1084_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _0627_ _0511_ _0744_ _0606_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3212_ _0205_ net71 u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2912__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _0139_ net74 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3074_ _0071_ net113 u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_SE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2025_ u_cpu.raddr\[1\] _0249_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1969__C _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2927_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _0229_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2858_ _0482_ _0529_ _0660_ _0689_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2356__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2789_ _1134_ _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1809_ _1218_ u_cpu.cpu.genblk3.csr.mcause31 _1248_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2903__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2595__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[19\] u_arbiter.i_wb_cpu_rdt\[16\] net128 u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ net14 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1570__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2681__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2712_ _0826_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2586__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2643_ _0455_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3228__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2338__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2574_ _0725_ _0726_ _0728_ _1382_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2338__B2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2889__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1561__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[52\]_CLK net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3126_ _0123_ net105 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2510__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[67\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3057_ _0054_ net89 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2008_ _0234_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2390__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2577__A1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2604__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__B2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2568__B2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2568__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ _0227_ u_arbiter.i_wb_cpu_rdt\[13\] _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_38_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2559__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0755_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2557_ _0571_ _0712_ _0649_ _0630_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2488_ _0490_ _0646_ _0649_ _0548_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3109_ _0106_ net79 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__B2 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2798__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2262__A3 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2970__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2005__A3 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _1214_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2261__I0 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout110_I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ u_cpu.cpu.decode.op21 _0486_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ _0425_ _0427_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2273_ _0227_ u_arbiter.i_wb_cpu_rdt\[0\] _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_42_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2229__B1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout23_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[20\]_SE net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__B _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1988_ u_cpu.cpu.immdec.imm11_7\[1\] _1398_ _1399_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2609_ u_cpu.cpu.immdec.imm19_12_20\[3\] _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2180__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2511__C _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2960_ _1002_ _1259_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2891_ net8 u_arbiter.o_wb_cpu_adr\[1\] _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[43\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1911_ _1335_ _1345_ _1346_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1842_ _1276_ _1280_ _1283_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1985__A2 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2934__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ u_cpu.cpu.bufreg2.i_cnt_done _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3236__D u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2325_ _0416_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2256_ _1091_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2187_ u_arbiter.i_wb_cpu_rdt\[15\] _0369_ _0370_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1988__B _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2870__B1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1900__A2 u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1664__A1 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1967__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1917__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1719__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[49\] u_scanchain_local.module_data_in\[48\] net135 u_arbiter.o_wb_cpu_adr\[11\]
+ net19 u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2392__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2144__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3153__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2110_ _0316_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3090_ _0087_ net51 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2041_ _0264_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__C _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2943_ _0987_ _0983_ _0991_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1958__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2080__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2874_ u_cpu.cpu.immdec.imm11_7\[2\] _0925_ _0945_ _0591_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ u_cpu.cpu.decode.co_ebreak _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1756_ u_arbiter.i_wb_cpu_dbus_adr\[29\] _1190_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ u_arbiter.i_wb_cpu_dbus_adr\[13\] _1143_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout90_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2308_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2239_ _1090_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2843__B1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2607__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2997__I1 u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3176__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2374__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2126__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2677__A3 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1885__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2517__B _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2062__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2590_ _0742_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3211_ _0204_ net70 u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3142_ _0014_ net75 u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3073_ _0070_ net112 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_cpu.rf_ram.RAM0_CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _0251_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2146__C _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3199__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2926_ _0978_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2053__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2857_ _0689_ _0429_ _0442_ _0498_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2788_ _0872_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1739_ u_arbiter.i_wb_cpu_dbus_adr\[25\] _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2903__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2044__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2595__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2347__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.output_buffers\[3\]_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2807__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2283__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2761__I _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0838_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2586__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2642_ _0413_ _0490_ _0502_ _0788_ _0574_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2573_ _0727_ _0726_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2338__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2001__I _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2897__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3125_ _0122_ net103 u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3056_ _0053_ net91 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1864__A4 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout53_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2007_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0236_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2274__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2026__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2909_ _0969_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2265__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2568__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2514__C _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[31\] u_arbiter.i_wb_cpu_rdt\[28\] net143 u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ net28 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2256__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2491__I _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2625_ _1237_ _0752_ _0773_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3237__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2192__B1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2556_ u_arbiter.i_wb_cpu_rdt\[29\] u_arbiter.i_wb_cpu_rdt\[13\] _0592_ _0712_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2487_ _0619_ _0528_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3108_ _0105_ net64 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3039_ _0036_ net72 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2247__A1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2798__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2970__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2486__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2238__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[51\]_CLK net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2410__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[66\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2961__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1655__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout103_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ _1268_ _0515_ _0578_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2687__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2341_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2272_ _1091_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_42_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2229__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[19\]_CLK net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout16_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _1392_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2608_ _0757_ _0752_ _0758_ _0559_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2539_ _0228_ u_arbiter.i_wb_cpu_rdt\[28\] _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2468__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2468__B2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[4\]_D u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3082__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1910_ _1331_ u_cpu.rf_ram_if.rdata1\[6\] _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2890_ _0723_ _0958_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ u_cpu.cpu.state.init_done _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1985__A3 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1772_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2324_ _0495_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2255_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2186_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _0375_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1988__C _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2870__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2622__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1664__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0262_ u_cpu.rf_ram.i_waddr\[1\] _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_u_scanchain_local.scan_flop\[10\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2764__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2852__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__C _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2942_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _1397_ _0982_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2080__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2873_ _0703_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1824_ _1263_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1755_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1686_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _1145_ _1142_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout83_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2307_ _0454_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2238_ _0411_ _0412_ _0413_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_39_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2169_ _0367_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2843__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_D u_arbiter.i_wb_cpu_rdt\[25\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__B _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2359__B1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1582__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2685__I1 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[19\]_D u_arbiter.i_wb_cpu_rdt\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[61\] u_scanchain_local.module_data_in\[60\] net141 u_arbiter.o_wb_cpu_adr\[23\]
+ net26 u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_16_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3120__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1573__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3210_ _0203_ net70 u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3141_ _0138_ net75 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3072_ _0069_ net112 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _0232_ _0245_ _0249_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_78_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2589__B1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2925_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0973_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2053__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2856_ _0630_ _0928_ _0552_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1807_ _1246_ _1247_ _1249_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_30_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2787_ _0886_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1738_ _1102_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[56\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1669_ _1135_ _1128_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3143__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2201__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout133_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _0833_
+ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1794__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2641_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_rdt\[1\] _0592_ _0788_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2572_ u_cpu.cpu.immdec.imm31 _1223_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2897__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3016__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3124_ _0121_ net103 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ _0052_ net89 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2006_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _0235_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2274__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout46_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2908_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _0967_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2577__A3 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2839_ _1397_ _1050_ _1229_ _1291_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2265__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2017__A2 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3039__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[24\] u_arbiter.i_wb_cpu_rdt\[21\] net131 u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ net16 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3189__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3080__D _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1700__A1 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2500__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ u_cpu.cpu.immdec.imm19_12_20\[5\] _0479_ _0771_ _0772_ _0755_ _0773_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2192__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2192__B2 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2555_ _0709_ _0469_ _0620_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2486_ _0543_ _0596_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3107_ _0104_ net63 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3038_ _0035_ net74 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2247__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1749__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2410__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2340_ _0230_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2271_ _0447_ _0441_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2477__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2229__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1988__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3204__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _1317_ _1215_ _1318_ _1309_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_120_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ u_cpu.cpu.immdec.imm19_12_20\[3\] _0509_ _0755_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2538_ _1095_ u_arbiter.i_wb_cpu_rdt\[12\] _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2469_ _1051_ _0591_ _0634_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2468__A2 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1979__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2951__I0 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1903__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ u_cpu.cpu.state.stage_two_req _1281_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2395__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ _1215_ u_cpu.cpu.bufreg.i_sh_signed _1048_ _1041_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_129_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2254_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2185_ _0378_ _0379_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_SE net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2870__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1969_ _1385_ _1270_ _1306_ _1372_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2386__A1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[7] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2377__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[18\]_CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2852__A2 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2941_ _1275_ _1372_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2604__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2872_ _0454_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2368__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1823_ _1264_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1754_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _1195_ _1196_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ _1145_ _1142_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1591__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout76_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2306_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2237_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0410_
+ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2168_ u_arbiter.i_wb_cpu_rdt\[10\] _0324_ _0326_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _0350_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2099_ _0282_ _1286_ _0035_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2690__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2359__A1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2359__B2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1582__A2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3072__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[54\] u_scanchain_local.module_data_in\[53\] net139 u_arbiter.o_wb_cpu_adr\[16\]
+ net23 u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2522__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3140_ _0137_ net112 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3071_ _0068_ net112 u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ u_cpu.raddr\[0\] _0247_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2589__B2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _0977_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2855_ _0461_ _0737_ _0777_ _0927_ _0517_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1806_ u_cpu.cpu.decode.op26 _1053_ _1049_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_121_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2786_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _0885_ _0880_ _1134_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1737_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1668_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ _1058_ _1077_ _1062_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2044__A3 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2201__B1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2752__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2504__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2807__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2544__B _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1794__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2640_ _0774_ _0785_ _0786_ _0787_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2571_ _1374_ _0297_ _1380_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3123_ _0120_ net98 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3054_ _0051_ net89 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2005_ u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[3\] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ net35 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_23_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout39_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[23\]_SE net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2907_ _0968_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ u_cpu.cpu.ctrl.i_jump _1294_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2769_ _1096_ _0870_ _0873_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[30\]_SI u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3110__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2973__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__A2 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[17\] u_arbiter.i_wb_cpu_rdt\[14\] net129 u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ net13 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1700__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2264__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ _0529_ _0504_ _0532_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2177__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2554_ _0423_ _0560_ _0611_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2192__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2485_ _0525_ _0599_ _0595_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3106_ _0103_ net63 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3037_ _0034_ net76 u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2955__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2168__C1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2183__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[69\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A1 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2238__A3 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2270_ _0226_ u_arbiter.i_wb_cpu_rdt\[14\] _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1985_ u_cpu.cpu.immdec.imm11_7\[4\] u_cpu.cpu.immdec.imm11_7\[3\] u_cpu.cpu.immdec.imm11_7\[2\]
+ u_cpu.cpu.immdec.imm11_7\[0\] _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_105_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ u_cpu.cpu.immdec.imm19_12_20\[2\] _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2165__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2537_ _0693_ _0694_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2468_ _0580_ _0608_ _0633_ _0606_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2399_ _0553_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3029__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1600__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3179__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1903__A2 u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2864__B1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1770_ u_arbiter.i_wb_cpu_dbus_we _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2395__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2322_ _0432_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2253_ _0410_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2184_ u_arbiter.i_wb_cpu_rdt\[14\] _0369_ _0370_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout21_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1968_ _1317_ _1380_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2386__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1899_ _1332_ _1337_ _1338_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1897__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2697__I0 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[6] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2129__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2598__I _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1888__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2301__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2065__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2940_ _0984_ _0983_ _0989_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2871_ _0549_ _0443_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1812__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__I _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1822_ u_cpu.cpu.decode.opcode\[0\] _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2368__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1753_ _1139_ _1200_ _1201_ u_arbiter.o_wb_cpu_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ _1124_ _1146_ _1148_ u_arbiter.o_wb_cpu_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2305_ _0434_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout69_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2236_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] _0410_
+ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ _0365_ _0366_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2098_ _0296_ _0309_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2056__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2359__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3217__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2295__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[47\] u_scanchain_local.module_data_in\[46\] net135 u_arbiter.o_wb_cpu_adr\[9\]
+ net19 u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3070_ _0067_ net117 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2021_ u_cpu.raddr\[0\] _0247_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2589__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2923_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _0973_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2854_ _0686_ _0626_ _0520_ _0481_ _0737_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1805_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2785_ _0868_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ _1185_ _1183_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1667_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1598_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ _0399_ _0361_ _0401_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3199_ _0192_ net82 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2277__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[17\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2201__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2752__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__A2 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2440__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2440__B2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1955__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout119_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ u_cpu.cpu.immdec.imm19_12_20\[0\] _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3122_ _0119_ net98 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3053_ _0050_ net89 u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2004_ _1282_ _0233_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3062__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2906_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2837_ u_cpu.cpu.ctrl.i_jump _1316_ _1050_ _1078_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2768_ _0875_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1719_ u_arbiter.i_wb_cpu_dbus_adr\[21\] _1147_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2699_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _0827_
+ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2498__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2422__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2380__B _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2489__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2555__B _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3085__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2264__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2964__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2622_ _0735_ _0765_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2177__B1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2553_ _0412_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2484_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _1093_ _0646_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3105_ _0102_ net63 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3036_ _0033_ net76 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_GWEN _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2652__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2404__B2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1809__B _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2168__B1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2359__C _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2891__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A2 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2238__A4 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2643__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[7\]_D u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[13\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2634__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1984_ _1078_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.out_flop_CLKN net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2304__I _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3100__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2605_ _0754_ _0752_ _0756_ _0551_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout99_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2536_ u_cpu.cpu.immdec.imm30_25\[2\] _0678_ _0679_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _0690_ _0580_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_2467_ _0629_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2398_ _0422_ _0518_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2873__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3019_ _0006_ net47 u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2625__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[36\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2864__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2864__B2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3123__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1963__I u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout101_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2321_ _0441_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _0425_ _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2183_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _0375_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2855__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2235__S _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout14_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1379_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2034__I _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2791__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1898_ _1335_ u_cpu.rf_ram_if.rdata1\[2\] _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2519_ _0570_ _0677_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1897__A2 u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1649__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2697__I1 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2637__C _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3146__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_WEN[5] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1585__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1888__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ u_cpu.cpu.immdec.imm11_7\[3\] _0479_ _0606_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ u_cpu.cpu.decode.opcode\[2\] _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2222__C1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1752_ u_arbiter.i_wb_cpu_dbus_adr\[28\] _1190_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1683_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3019__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2304_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2235_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0410_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2166_ u_arbiter.i_wb_cpu_rdt\[9\] _0343_ _0352_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2029__I _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ _0297_ _0308_ _0028_ _1373_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2999_ u_cpu.rf_ram_if.wdata0_r\[5\] u_cpu.rf_ram_if.wdata1_r\[5\] _1020_ _1028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3005__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_cpu.rf_ram.RAM0 u_cpu.rf_ram.RAM0/A[0] u_cpu.rf_ram.RAM0/A[1] u_cpu.rf_ram.RAM0/A[2]
+ u_cpu.rf_ram.RAM0/A[3] u_cpu.rf_ram.RAM0/A[4] u_cpu.rf_ram.RAM0/A[5] u_cpu.rf_ram.RAM0/A[6]
+ u_cpu.rf_ram.RAM0/A[7] u_cpu.rf_ram.RAM0/CEN u_cpu.rf_ram.RAM0/CLK u_cpu.rf_ram.RAM0/D[0]
+ u_cpu.rf_ram.RAM0/D[1] u_cpu.rf_ram.RAM0/D[2] u_cpu.rf_ram.RAM0/D[3] u_cpu.rf_ram.RAM0/D[4]
+ u_cpu.rf_ram.RAM0/D[5] u_cpu.rf_ram.RAM0/D[6] u_cpu.rf_ram.RAM0/D[7] u_cpu.rf_ram.RAM0/GWEN
+ u_cpu.rf_ram.RAM0/Q[0] u_cpu.rf_ram.RAM0/Q[1] u_cpu.rf_ram.RAM0/Q[2] u_cpu.rf_ram.RAM0/Q[3]
+ u_cpu.rf_ram.RAM0/Q[4] u_cpu.rf_ram.RAM0/Q[5] u_cpu.rf_ram.RAM0/Q[6] u_cpu.rf_ram.RAM0/Q[7]
+ u_cpu.rf_ram.RAM0/WEN[0] u_cpu.rf_ram.RAM0/WEN[1] u_cpu.rf_ram.RAM0/WEN[2] u_cpu.rf_ram.RAM0/WEN[3]
+ u_cpu.rf_ram.RAM0/WEN[4] u_cpu.rf_ram.RAM0/WEN[5] u_cpu.rf_ram.RAM0/WEN[6] u_cpu.rf_ram.RAM0/WEN[7]
+ vdd vss gf180mcu_fd_ip_sram__sram256x8m8wm1
XFILLER_33_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2020_ _0246_ _0247_ _0248_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2922_ _0976_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2853_ _1219_ _0925_ _0926_ _0745_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1804_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2784_ _0884_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ _1172_ _1186_ _1187_ u_arbiter.o_wb_cpu_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ u_arbiter.i_wb_cpu_dbus_adr\[10\] _1103_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1597_ u_cpu.cpu.immdec.imm19_12_20\[5\] _1038_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout81_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ u_arbiter.i_wb_cpu_rdt\[26\] _0328_ _0400_ u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3198_ _0191_ net82 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2149_ _0351_ _0353_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1788__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2201__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1712__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2097__C _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A1 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2440__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3121_ _0118_ net98 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3052_ _0049_ net87 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2003_ _1298_ _1279_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3207__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2751__B _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2905_ _0229_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2836_ _0914_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2767_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0870_ _0873_ _1096_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2042__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1718_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2698_ _0831_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1649_ u_arbiter.i_wb_cpu_dbus_adr\[6\] _1115_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2498__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2422__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2186__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2489__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2110__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2571__B _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2177__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2621_ _0766_ _0739_ _0769_ _0483_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2177__B2 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ _0512_ _0696_ _0705_ _0708_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2797__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ _0643_ _0638_ _0645_ _0607_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[16\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3104_ _0101_ net49 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3035_ _0032_ net76 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout44_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2652__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2404__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2168__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2819_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _0899_ _0901_ _1185_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[22\] u_arbiter.i_wb_cpu_rdt\[19\] net131 u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ net16 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_61_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2331__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2634__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1983_ _1065_ _1396_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2604_ u_cpu.cpu.immdec.imm19_12_20\[2\] _0509_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2535_ _0685_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2466_ _0630_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2397_ _0445_ _0467_ _0498_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2322__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3018_ _0005_ net47 u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2990__I _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2389__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2431__S _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout151 net4 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2864__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2386__B _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2927__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2320_ _0493_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2552__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2182_ _0376_ _0377_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2855__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2315__I _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1966_ _1232_ _1381_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1897_ _1333_ u_cpu.rf_ram.rdata\[2\] _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3098__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1594__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[9\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0538_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2449_ _0531_ _0613_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_WEN[4] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2231__B1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2534__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2534__B2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2837__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[10\]_SI u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3240__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1820_ _1041_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2222__B1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2222__C2 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1751_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1576__A2 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1682_ _1102_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2303_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ u_arbiter.i_wb_cpu_rdt\[11\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _0361_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2096_ _1241_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[26\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3005__A2 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ _1027_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1949_ _1361_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_33_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2516__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3113__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2755__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1730__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0973_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2852_ u_cpu.cpu.immdec.imm11_7\[1\] _0644_ _0924_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2783_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _0878_ _0880_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1803_ u_cpu.cpu.decode.op22 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1734_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _1147_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1665_ _1124_ _1131_ _1132_ u_arbiter.o_wb_cpu_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1596_ _1038_ _1050_ _1073_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _1282_ _0243_ _0314_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3197_ _0190_ net82 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2148_ u_arbiter.i_wb_cpu_rdt\[4\] _0343_ _0352_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2079_ _0292_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2704__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1828__B u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1960__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2673__B1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3009__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2976__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1779__A2 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2189__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[52\] u_scanchain_local.module_data_in\[51\] net136 u_arbiter.o_wb_cpu_adr\[14\]
+ net19 u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3159__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3120_ _0117_ net96 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1703__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3051_ _0048_ net91 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ _1077_ u_cpu.cpu.state.stage_two_req _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_97_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2967__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0966_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2751__C _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2835_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _0869_ _0872_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2766_ _0874_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1717_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _1167_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2697_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _0827_
+ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1648_ _1087_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1942__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ u_cpu.cpu.genblk3.csr.o_new_irq _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3249_ _0222_ net40 u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2670__A3 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2258__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2958__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2233__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2186__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2389__B _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1697__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2620_ _0735_ _0737_ _0767_ _0768_ _0597_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2177__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1982__I _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ u_cpu.cpu.immdec.imm30_25\[3\] _0706_ _0707_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2482_ u_cpu.cpu.immdec.imm24_20\[3\] _0636_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2724__I1 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1688__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3103_ _0100_ net63 u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3034_ _0031_ net74 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2101__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2318__I _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout37_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2254__S _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2818_ _0904_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2168__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2749_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2988__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1892__I _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2002__B _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1679__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2715__I1 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2656__C _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2651__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__A2 u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[15\] u_arbiter.i_wb_cpu_rdt\[12\] net129 u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ net13 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_42_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2331__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.input_buf_clk net1 u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1982_ _1370_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2603_ _0750_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2534_ _0687_ _0688_ _0691_ _0587_ _0673_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2465_ _0560_ _0543_ _0448_ _0608_ _0548_ _0627_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_2396_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _1094_ _0565_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2858__B1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2322__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3017_ _0004_ net41 u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1833__A1 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2389__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1836__B _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2010__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[62\]_CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2561__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout130 net133 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout141 net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2077__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1824__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[15\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2927__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _0420_ u_arbiter.i_wb_cpu_rdt\[1\] _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2181_ u_arbiter.i_wb_cpu_rdt\[13\] _0369_ _0370_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2068__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1815__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1815__B2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1965_ _1328_ _1265_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1896_ _1332_ _1334_ _1336_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2517_ _0297_ _0676_ _1369_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2448_ _0598_ _0613_ _0458_ _0494_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2379_ _0474_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_WEN[3] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2442__S _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2231__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3042__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2231__B2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_scanchain_local.scan_flop\[8\] u_arbiter.i_wb_cpu_rdt\[5\] net132 u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ net15 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_102_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2222__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1750_ _1195_ _1196_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2151__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1681_ _1145_ _1142_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2525__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2302_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2289__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2233_ u_cpu.cpu.genblk1.align.ctrl_misal _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2164_ _0364_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2095_ _0302_ _0304_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3065__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2997_ _1026_ u_cpu.rf_ram.i_wdata\[4\] _1022_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1948_ _1368_ u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_102_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1879_ _1321_ u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.bufreg.lsb\[1\]
+ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2010__B u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2452__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2204__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2755__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3088__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2574__C _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2920_ _0975_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[8\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2851_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2782_ _0883_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1802_ u_cpu.cpu.state.o_cnt_r\[3\] _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ _1185_ _1183_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2746__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1664_ u_arbiter.i_wb_cpu_dbus_adr\[9\] _1115_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1595_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _1054_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2216_ u_arbiter.i_wb_cpu_dbus_dat\[27\] _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3196_ _0189_ net82 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout67_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2147_ _0325_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2078_ _1085_ u_cpu.cpu.state.o_cnt_r\[2\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1844__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3230__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2673__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2673__B2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2189__C2 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2189__B1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[30\]_D u_arbiter.i_wb_cpu_rdt\[27\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[45\] u_scanchain_local.module_data_in\[44\] net138 u_arbiter.o_wb_cpu_adr\[7\]
+ net22 u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_103_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[16\]_SE net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3050_ _0047_ net88 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ _0230_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2664__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2416__A1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2903_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _0961_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[23\]_SI u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2834_ _0913_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_D u_arbiter.i_wb_cpu_rdt\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2765_ _1084_ _0870_ _0873_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1716_ _1105_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2696_ _0830_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1647_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _1112_ _1113_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1578_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3248_ _0221_ net40 u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3179_ _0173_ net50 u_cpu.rf_ram.i_waddr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2655__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2715__S _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2258__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[12\]_D u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[39\]_SE net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3126__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2424__I _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout117_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2550_ _0532_ _0677_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ _0478_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2885__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3102_ _0099_ net63 u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3033_ _0030_ net74 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2637__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1860__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2817_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _0899_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2748_ _0826_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2679_ u_cpu.cpu.alu.cmp_r _1370_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2876__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[69\]_SI u_arbiter.o_wb_cpu_adr\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2628__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3149__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2651__I1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2619__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ _1394_ _1395_ _1393_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2602_ u_cpu.cpu.immdec.imm19_12_20\[1\] _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2533_ _0689_ _0610_ _0690_ _0660_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2103__B _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2464_ _0503_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2858__B2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2395_ _1059_ _0515_ _0564_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3016_ _0003_ net41 u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2492__C _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2948__B _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2561__A3 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout120 net121 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2849__A1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout142 net150 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_130_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _1263_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1895_ _1335_ u_cpu.rf_ram_if.rdata1\[1\] _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout97_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ _1372_ _1374_ _1215_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2447_ _0462_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2378_ _0423_ _0540_ _0546_ _0517_ _0548_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_42_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_WEN[2] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3008__A1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2231__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2767__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2222__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1680_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2301_ net8 _1086_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2232_ _0407_ _0352_ _0409_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2163_ u_arbiter.i_wb_cpu_rdt\[8\] _0324_ _0326_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _0350_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_22_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2094_ _1296_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[61\]_CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout12_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ u_cpu.rf_ram_if.wdata0_r\[4\] u_cpu.rf_ram_if.wdata1_r\[4\] _1020_ _1026_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1947_ u_cpu.rf_ram_if.rtrig0 _1066_ _1362_ u_cpu.rf_ram.i_waddr\[7\] _1368_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1878_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2516__A3 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2498__B _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[14\]_CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[29\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2961__B _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2204__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1715__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2140__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2855__C _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2850_ _0231_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1801_ _1244_ _1239_ _1241_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2781_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _0878_ _0880_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1732_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _1128_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1594_ u_cpu.cpu.immdec.imm24_20\[1\] _1065_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _0398_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3032__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3195_ _0188_ net84 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2146_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0320_ _0348_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ _0281_ _1311_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2337__I _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3182__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2434__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2979_ _1015_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2800__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1844__C _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2956__B _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2122__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2673__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2189__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2189__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[38\] u_scanchain_local.module_data_in\[37\] net132 u_arbiter.o_wb_cpu_adr\[0\]
+ net15 u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3055__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2361__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2000_ _0228_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0229_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2664__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2902_ _0965_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1996__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2833_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0869_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2764_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1715_ _1124_ _1170_ _1171_ u_arbiter.o_wb_cpu_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2695_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _0827_ _0830_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1646_ _1112_ _1113_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1577_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3247_ _0220_ net39 u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3178_ _0172_ net102 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2655__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2129_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _1321_ net35 _0317_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2407__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2591__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3078__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__B2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[7\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A3 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2906__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1909__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2582__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2480_ u_cpu.cpu.immdec.imm24_20\[2\] _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3101_ _0098_ net44 u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2885__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3032_ _0029_ net76 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2637__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2816_ _0903_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ u_cpu.cpu.bufreg.i_sh_signed _1400_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2678_ _0818_ _0819_ _0820_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2573__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1629_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2876__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[0\]_SE net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2564__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2316__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2867__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2619__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1980_ _1314_ _1315_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ _0725_ _0752_ _0753_ _0578_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2532_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _0592_ _0690_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2555__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2463_ _0612_ _0625_ _0628_ _0492_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2858__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2394_ _0474_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3015_ _0002_ net41 u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[29\]_SE net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout42_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1833__A3 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1597__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2546__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout110 net111 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3116__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2849__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout143 net146 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout132 net133 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2255__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2537__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[20\] u_arbiter.i_wb_cpu_rdt\[17\] net129 u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ net13 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1760__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ u_cpu.cpu.decode.opcode\[1\] _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _1331_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3139__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2515_ _0672_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2446_ _0609_ _0611_ _0470_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2377_ _0450_ _0452_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[1] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1806__A3 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1990__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2519__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2914__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[68\] u_scanchain_local.module_data_in\[67\] net147 u_arbiter.o_wb_cpu_adr\[30\]
+ net30 u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2758__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2930__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2300_ _0420_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2231_ u_arbiter.i_wb_cpu_rdt\[31\] _0321_ _0405_ _1230_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2162_ _0362_ _0363_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2093_ u_cpu.cpu.alu.cmp_r _1306_ _0303_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2749__A1 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2995_ _1025_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1946_ _1071_ _1362_ _1367_ u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1877_ _1241_ u_cpu.cpu.mem_bytecnt\[0\] u_cpu.cpu.mem_bytecnt\[1\] _1320_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1972__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2429_ _0549_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2437__B1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2443__I _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2780_ _0882_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _1103_ _1181_ _1183_ _1184_ u_arbiter.o_wb_cpu_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1662_ _1124_ _1129_ _1130_ u_arbiter.o_wb_cpu_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1593_ _1070_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3194_ _0187_ net90 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2214_ u_arbiter.i_wb_cpu_rdt\[25\] _0372_ _0359_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _0373_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2145_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2076_ _0291_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2353__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2978_ _1333_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram_if.rtrig0 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_33_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2198__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2442__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1929_ _1356_ u_cpu.rf_ram_if.rtrig1 _1038_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_33_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2528__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1881__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2681__I0 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2189__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1607__I u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[60\]_CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2361__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1872__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2901_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _0961_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1624__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2672__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[62\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ _0912_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2763_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[13\]_CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1714_ u_arbiter.i_wb_cpu_dbus_adr\[20\] _1147_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2694_ _0829_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1645_ _1106_ _1114_ _1116_ u_arbiter.o_wb_cpu_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[28\]_CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1576_ u_cpu.cpu.decode.co_ebreak _1052_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2352__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout72_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3246_ _0219_ net37 u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2104__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ _0171_ net112 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2128_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _0317_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2059_ u_cpu.cpu.mem_bytecnt\[0\] _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2591__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1854__A1 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2803__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[50\] u_scanchain_local.module_data_in\[49\] net135 u_arbiter.o_wb_cpu_adr\[12\]
+ net20 u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1909__A2 u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3172__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3100_ _0097_ net44 u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3031_ _0028_ net72 u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1845__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1800__I _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _0899_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2746_ _1384_ _1387_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2022__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2677_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1628_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2325__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1559_ u_cpu.cpu.bufreg.lsb\[0\] _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3229_ _0212_ net55 u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1836__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3045__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2013__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3195__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2564__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2917__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2252__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout122_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2004__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ u_cpu.cpu.immdec.imm19_12_20\[1\] _0509_ _0751_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2531_ _0418_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2555__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2462_ _0438_ _0626_ _0520_ _0627_ _0428_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2393_ _0560_ _0453_ _0562_ _0517_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3014_ _0001_ net47 u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3068__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1833__A4 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[6\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2546__A2 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2729_ _0848_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout122 net123 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout111 net122 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout100 net101 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout144 net146 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout133 net134 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2737__S _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2980__B _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1615__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[13\] u_arbiter.i_wb_cpu_rdt\[10\] net128 u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ net12 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3210__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2225__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1962_ u_cpu.cpu.bufreg.c_r _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1893_ _1333_ u_cpu.rf_ram.rdata\[1\] _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2514_ _0423_ _0527_ _0582_ _0491_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2445_ _0467_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2161__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2376_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_WEN[0] _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2519__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2959__C _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3233__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[0\]_D net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2455__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_u_scanchain_local.scan_flop\[19\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _0407_ _0361_ _0408_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.out_flop_D u_scanchain_local.module_data_in\[69\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2161_ u_arbiter.i_wb_cpu_rdt\[7\] _0343_ _0352_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2092_ _0299_ _0301_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2176__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2446__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2994_ _1024_ u_cpu.rf_ram.i_wdata\[3\] _1022_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2125__B _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1945_ u_cpu.rf_ram.i_waddr\[6\] _1358_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ u_cpu.cpu.mem_if.signbit _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2428_ _0567_ _0583_ _0470_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2359_ _0527_ _0529_ _0455_ _0531_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2437__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2437__B2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[6\] u_arbiter.i_wb_cpu_rdt\[3\] net126 u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ net9 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2676__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2925__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[33\]_D u_arbiter.i_wb_cpu_rdt\[30\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1730_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _1123_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ u_arbiter.i_wb_cpu_dbus_adr\[8\] _1115_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1592_ u_cpu.cpu.immdec.imm19_12_20\[8\] _1068_ _1069_ u_cpu.cpu.immdec.imm24_20\[4\]
+ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3193_ _0186_ net84 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2213_ _0396_ _0397_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2667__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2144_ _0243_ _0315_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2075_ _0279_ _1290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_74_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[24\]_D u_arbiter.i_wb_cpu_rdt\[21\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2977_ _0245_ _1014_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2442__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1928_ u_cpu.rf_ram_if.o_wen_req _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1859_ _1299_ _1300_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2809__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[15\]_D u_arbiter.i_wb_cpu_rdt\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A1 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _0964_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2831_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _0906_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2762_ net2 _1393_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _1167_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2693_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _0827_ _0829_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1644_ u_arbiter.i_wb_cpu_dbus_adr\[5\] _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1575_ _1053_ _1049_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2352__A3 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3245_ _0218_ net37 u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3176_ _0170_ net118 u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout65_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ _0334_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1863__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2058_ _0272_ _0276_ _0277_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2364__I _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2879__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1618__I _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[43\] u_scanchain_local.module_data_in\[42\] net137 u_arbiter.o_wb_cpu_adr\[5\]
+ net21 u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1790__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3030_ _0012_ net45 u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1845__A2 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2270__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ _0902_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _1384_ _1387_ _1400_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ _0273_ _1400_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1627_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1558_ _1038_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3228_ u_cpu.rf_ram_if.rtrig0 net48 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3159_ _0153_ net96 u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2013__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2043__B _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1772__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__B _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1827__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[27\]_CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2004__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout115_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _0482_ _0626_ _0428_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2461_ _0414_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2563__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2392_ _0435_ _0464_ _0554_ _0561_ _0553_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2179__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3013_ _0000_ net47 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1818__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout28_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _0845_
+ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2659_ _0774_ _0802_ _0803_ _0804_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xfanout112 net114 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout101 net102 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout145 net149 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout134 net151 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3012__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2482__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3162__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1993__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2170__A1 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2225__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1961_ _1302_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _1226_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2513_ _0506_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2444_ _0465_ _0496_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3035__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2375_ _0493_ _0501_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2161__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1716__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1966__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3058__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2930__A3 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2160_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2091_ _1236_ _1244_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2446__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2993_ u_cpu.rf_ram_if.wdata0_r\[3\] u_cpu.rf_ram_if.wdata1_r\[3\] _1020_ _1024_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1944_ _1070_ _1361_ _1366_ u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_33_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1875_ _1263_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout95_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2427_ _0574_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ _0478_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2289_ _1091_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3200__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2373__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2676__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1939__A1 u_cpu.rf_ram.i_waddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2600__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1660_ _1127_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1591_ u_cpu.cpu.immdec.imm19_12_20\[7\] _1068_ _1069_ u_cpu.cpu.immdec.imm24_20\[3\]
+ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2116__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3192_ _0185_ net90 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2212_ u_arbiter.i_wb_cpu_rdt\[24\] _0386_ _0357_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2143_ _0320_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2074_ _0287_ _0290_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3223__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout10_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2976_ _0232_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1927_ _1347_ _1345_ _1355_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1858_ _1284_ _1283_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1789_ _1217_ _1231_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2298__S _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[3\]_SE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2594__B2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2649__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3246__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ _0911_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout145_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2761_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2692_ _0828_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1712_ _1154_ _1167_ _1168_ _1169_ u_arbiter.o_wb_cpu_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2585__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1643_ _1102_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1574_ _1041_ u_cpu.cpu.decode.opcode\[2\] _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2888__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3244_ _0217_ net36 u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3175_ _0169_ net118 u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2126_ u_arbiter.i_wb_cpu_rdt\[1\] _0328_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout58_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2057_ _1246_ u_cpu.cpu.state.o_cnt\[2\] _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2959_ _0273_ _1261_ _1002_ _1251_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_124_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2328__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3119__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2879__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2803__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2031__A3 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[36\] u_scanchain_local.module_data_in\[35\] net145 u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ net27 u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__A3 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2813_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _0899_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2558__B2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2558__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2744_ _0856_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2675_ u_cpu.cpu.genblk3.csr.timer_irq_r _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1626_ _1085_ u_cpu.cpu.state.ibus_cyc _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1557_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_28_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3227_ _0211_ net71 u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3158_ _0152_ net96 u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2109_ _1321_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1836__A3 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3089_ _0086_ net51 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2549__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1882__C _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3091__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2260__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1763__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2460_ _0458_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2563__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2391_ _0536_ _0531_ _0524_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3012_ _0022_ net54 u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2195__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _0847_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2658_ u_cpu.cpu.immdec.imm19_12_20\[7\] _0751_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1609_ _1085_ u_cpu.cpu.state.ibus_cyc _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfanout102 net111 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_2589_ _0445_ _0571_ _0660_ _0627_ _0575_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_43_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout146 net149 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout124 net5 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout135 net137 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2170__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1912__I _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _1377_ _1087_ u_arbiter.o_wb_cpu_we vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1891_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _0492_ _0670_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2443_ _0598_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2374_ _0438_ _0464_ _0541_ _0542_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_25_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2161__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2139__B _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout40_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[42\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[26\]_CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2049__B _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1888__B _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2090_ _0299_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_111_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[65\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2992_ _1023_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ u_cpu.rf_ram.i_waddr\[5\] _1358_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1874_ _1265_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1817__I _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2426_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _0592_ _0593_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout88_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3152__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2357_ _0228_ u_arbiter.i_wb_cpu_rdt\[5\] _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2288_ _0431_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1893__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2693__I0 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2383__I _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1884__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1636__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[66\] u_scanchain_local.module_data_in\[65\] net148 u_arbiter.o_wb_cpu_adr\[28\]
+ net31 u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2061__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1939__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3025__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3175__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1590_ _1067_ _1066_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_84_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2116__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3191_ _0184_ net84 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2211_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0352_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2142_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _0235_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2521__C1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1875__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2073_ _0279_ _1396_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2975_ _0225_ u_cpu.rf_ram_if.rcnt\[1\] _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1926_ u_cpu.rf_ram_if.rdata0\[7\] _1350_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1857_ _1212_ _1279_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1991__B _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1788_ _1232_ u_cpu.cpu.alu.add_cy_r _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2409_ _0511_ _0565_ _0569_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_44_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2291__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3198__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2043__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2288__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1857__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1609__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2282__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2760_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout138_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2691_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _0827_ _0828_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1711_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _1123_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2585__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1642_ _1112_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1573_ u_cpu.cpu.decode.op21 _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3243_ _0216_ net36 u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3174_ _0168_ net118 u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2125_ _0329_ _0331_ _0321_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2056_ _1246_ u_cpu.cpu.state.o_cnt\[2\] _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2273__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2958_ _1061_ _1254_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1909_ _1226_ u_cpu.rf_ram.rdata\[6\] _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2889_ u_cpu.cpu.bufreg.i_sh_signed _0480_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2328__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2879__A3 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2610__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1839__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2016__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2031__A4 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[29\] u_arbiter.i_wb_cpu_rdt\[26\] net133 u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ net16 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3213__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2007__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2812_ _0871_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2743_ u_arbiter.i_wb_cpu_dbus_adr\[30\] u_arbiter.i_wb_cpu_dbus_adr\[31\] _0851_
+ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2674_ _0480_ _0612_ _0815_ _0817_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1625_ _1087_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1825__I u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1556_ u_cpu.rf_ram_if.rcnt\[2\] _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout70_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3226_ _0210_ net45 u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3157_ _0151_ net97 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2108_ _0234_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3088_ _0085_ net50 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2039_ _0254_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3236__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2485__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2960__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2173__B1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2390_ _0493_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3011_ _0021_ net54 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3109__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2726_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _0845_
+ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2400__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ u_cpu.cpu.immdec.imm19_12_20\[8\] _0514_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1608_ net2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout103 net105 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2588_ _0489_ _0733_ _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout114 net117 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout147 net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout125 net127 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout136 net137 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3209_ _0202_ net58 u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2942__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[3\]_D u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2630__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1890_ u_cpu.rf_ram_if.rtrig1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout120_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2511_ _0609_ _0616_ _0620_ _0567_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_83_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2442_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _1093_ _0608_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2373_ _0524_ _0544_ _0448_ _0542_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2449__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout33_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3081__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__B _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2709_ _0837_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1888__C _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2860__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1966__A3 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A3 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[11\] u_arbiter.i_wb_cpu_rdt\[8\] net125 u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ net10 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_79_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2991_ _1021_ u_cpu.rf_ram.i_wdata\[2\] _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _1081_ _1361_ _1365_ u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1873_ _1314_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1957__A3 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3237__D u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2425_ _1093_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1590__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2356_ _1092_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2287_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1893__A2 u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1989__B _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2693__I1 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[27\]_D u_arbiter.i_wb_cpu_rdt\[24\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_cpu.rf_ram.RAM0_152 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[18\]_D u_arbiter.i_wb_cpu_rdt\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[59\] u_scanchain_local.module_data_in\[58\] net140 u_arbiter.o_wb_cpu_adr\[21\]
+ net23 u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2210_ _0394_ _0395_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3190_ _0183_ net84 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2521__B1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _0341_ _0343_ _0345_ _0346_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2685__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1875__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2072_ _0288_ _0245_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[10\]_CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2974_ _1012_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_u_scanchain_local.scan_flop\[25\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1925_ _1347_ _1343_ _1354_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1856_ _1058_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _1263_ _1298_ _1299_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ u_cpu.cpu.alu.i_rs1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1563__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2408_ _0570_ _0504_ _0573_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2339_ _0488_ _0508_ _0513_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2291__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2043__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[55\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[4\] u_arbiter.i_wb_cpu_rdt\[1\] net125 u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ net9 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_21_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3142__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1710_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _1164_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2690_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1641_ u_cpu.cpu.genblk1.align.ctrl_misal u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1572_ u_cpu.cpu.decode.op26 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3242_ _0215_ net71 u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input5_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3173_ _0167_ net109 u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2124_ net35 _0319_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1848__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2055_ _0275_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2273__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1986__C _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2957_ _0998_ _1000_ _1001_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1558__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1908_ _1332_ _1343_ _1344_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2888_ _0952_ _0925_ _0956_ _0957_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1839_ _1264_ _1046_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1784__A1 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3015__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2016__A2 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout150_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ _0900_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2742_ _0855_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2673_ u_cpu.cpu.immdec.imm31 _0509_ _0580_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1624_ _1098_ _1096_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3038__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1555_ u_cpu.rf_ram_if.rcnt\[0\] _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3225_ u_cpu.rf_ram_if.wtrig0 net48 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[3\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3156_ _0150_ net97 u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2107_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3087_ _0084_ net56 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2038_ u_cpu.raddr\[1\] _0261_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_19_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1757__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2485__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[41\] u_scanchain_local.module_data_in\[40\] net137 u_arbiter.o_wb_cpu_adr\[3\]
+ net21 u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2173__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3010_ _0020_ net54 u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0846_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2441__B _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2656_ _0484_ _0797_ _0801_ _0653_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_47_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1607_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout104 net105 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2587_ _0735_ _0737_ _0738_ _0740_ _0597_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout115 net116 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout126 net127 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout137 net142 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1911__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout148 net149 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3208_ _0201_ net58 u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3139_ _0136_ net118 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2219__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2702__I0 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2526__B _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2630__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0445_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2394__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ _1247_ _0591_ _0607_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2146__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2372_ _0436_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3226__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout26_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2708_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _0833_
+ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2639_ u_cpu.cpu.immdec.imm19_12_20\[5\] _0774_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2999__I0 u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2128__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2679__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2923__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3249__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2990_ _0254_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_128_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ u_cpu.rf_ram.i_waddr\[4\] _1358_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1872_ _1084_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2367__B2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _0538_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2914__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2355_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2286_ _0459_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2833__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2597__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1934__I _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3071__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2521__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2140_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _0337_ _0342_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2071_ u_cpu.rf_ram_if.rgnt _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2973_ _0279_ u_cpu.rf_ram_if.rreq_r _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2588__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1924_ u_cpu.rf_ram_if.rdata0\[6\] _1350_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1855_ _1058_ u_cpu.cpu.state.init_done _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ _1216_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2512__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2407_ _0445_ _0541_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2338_ _1374_ _0509_ _0435_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2269_ _1090_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2028__B1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2579__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3094__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1690__S _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2503__A1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1640_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1571_ u_cpu.cpu.decode.op21 _1044_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_119_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3241_ _0214_ net46 u_cpu.rf_ram_if.o_wen_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3172_ _0166_ net109 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2123_ _0316_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ _0272_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2956_ _1259_ _1000_ _0279_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1907_ _1331_ u_cpu.rf_ram_if.rdata1\[5\] _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2887_ u_cpu.cpu.immdec.imm30_25\[0\] _0486_ _0925_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1838_ _1045_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2981__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1784__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1769_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_SE net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput6 net6 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[24\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[39\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout143_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2810_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _0899_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2741_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[30\] _0851_
+ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2672_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _1095_ _0816_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.output_buffers\[3\] net31 u_scanchain_local.clk_out vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1623_ _1094_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_12_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ u_cpu.rf_ram_if.rcnt\[1\] _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2191__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3224_ u_cpu.cpu.o_wdata0 net46 u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
.ends

