// This is the unpowered netlist.
module serv_0 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_arbiter.o_wb_cpu_adr[0] ;
 wire \u_arbiter.o_wb_cpu_adr[10] ;
 wire \u_arbiter.o_wb_cpu_adr[11] ;
 wire \u_arbiter.o_wb_cpu_adr[12] ;
 wire \u_arbiter.o_wb_cpu_adr[13] ;
 wire \u_arbiter.o_wb_cpu_adr[14] ;
 wire \u_arbiter.o_wb_cpu_adr[15] ;
 wire \u_arbiter.o_wb_cpu_adr[16] ;
 wire \u_arbiter.o_wb_cpu_adr[17] ;
 wire \u_arbiter.o_wb_cpu_adr[18] ;
 wire \u_arbiter.o_wb_cpu_adr[19] ;
 wire \u_arbiter.o_wb_cpu_adr[1] ;
 wire \u_arbiter.o_wb_cpu_adr[20] ;
 wire \u_arbiter.o_wb_cpu_adr[21] ;
 wire \u_arbiter.o_wb_cpu_adr[22] ;
 wire \u_arbiter.o_wb_cpu_adr[23] ;
 wire \u_arbiter.o_wb_cpu_adr[24] ;
 wire \u_arbiter.o_wb_cpu_adr[25] ;
 wire \u_arbiter.o_wb_cpu_adr[26] ;
 wire \u_arbiter.o_wb_cpu_adr[27] ;
 wire \u_arbiter.o_wb_cpu_adr[28] ;
 wire \u_arbiter.o_wb_cpu_adr[29] ;
 wire \u_arbiter.o_wb_cpu_adr[2] ;
 wire \u_arbiter.o_wb_cpu_adr[30] ;
 wire \u_arbiter.o_wb_cpu_adr[31] ;
 wire \u_arbiter.o_wb_cpu_adr[3] ;
 wire \u_arbiter.o_wb_cpu_adr[4] ;
 wire \u_arbiter.o_wb_cpu_adr[5] ;
 wire \u_arbiter.o_wb_cpu_adr[6] ;
 wire \u_arbiter.o_wb_cpu_adr[7] ;
 wire \u_arbiter.o_wb_cpu_adr[8] ;
 wire \u_arbiter.o_wb_cpu_adr[9] ;
 wire \u_arbiter.o_wb_cpu_cyc ;
 wire \u_arbiter.o_wb_cpu_we ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.addr[0] ;
 wire \u_cpu.rf_ram.addr[1] ;
 wire \u_cpu.rf_ram.addr[2] ;
 wire \u_cpu.rf_ram.addr[3] ;
 wire \u_cpu.rf_ram.addr[4] ;
 wire \u_cpu.rf_ram.addr[5] ;
 wire \u_cpu.rf_ram.addr[6] ;
 wire \u_cpu.rf_ram.addr[7] ;
 wire \u_cpu.rf_ram.data[0] ;
 wire \u_cpu.rf_ram.data[1] ;
 wire \u_cpu.rf_ram.data[2] ;
 wire \u_cpu.rf_ram.data[3] ;
 wire \u_cpu.rf_ram.data[4] ;
 wire \u_cpu.rf_ram.data[5] ;
 wire \u_cpu.rf_ram.data[6] ;
 wire \u_cpu.rf_ram.data[7] ;
 wire \u_cpu.rf_ram.i_wdata[0] ;
 wire \u_cpu.rf_ram.i_wdata[1] ;
 wire \u_cpu.rf_ram.i_wdata[2] ;
 wire \u_cpu.rf_ram.i_wdata[3] ;
 wire \u_cpu.rf_ram.i_wdata[4] ;
 wire \u_cpu.rf_ram.i_wdata[5] ;
 wire \u_cpu.rf_ram.i_wdata[6] ;
 wire \u_cpu.rf_ram.i_wdata[7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.clk ;
 wire \u_scanchain_local.clk_out ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.data_out_i ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1357_ (.I(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1358_ (.I(\u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1359_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0849_),
    .A3(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1360_ (.I(_0851_),
    .ZN(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1361_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1362_ (.A1(_0852_),
    .A2(\u_cpu.cpu.bufreg.lsb[1] ),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1363_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1364_ (.I(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1365_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1366_ (.I(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1367_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1368_ (.I(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1369_ (.A1(_0856_),
    .A2(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1370_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1371_ (.A1(_0860_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1372_ (.A1(_0854_),
    .A2(\u_cpu.cpu.decode.op21 ),
    .A3(_0859_),
    .A4(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1373_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1374_ (.I(\u_cpu.cpu.decode.op21 ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1375_ (.A1(_0864_),
    .A2(\u_cpu.cpu.decode.op26 ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1376_ (.A1(_0854_),
    .A2(_0861_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1377_ (.A1(_0859_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1378_ (.A1(_0863_),
    .A2(_0865_),
    .B(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1379_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1380_ (.A1(_0855_),
    .A2(_0857_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1381_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_0870_),
    .A3(_0866_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1382_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1383_ (.A1(_0869_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1384_ (.A1(_0868_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1385_ (.A1(_0862_),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1386_ (.A1(_0851_),
    .A2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1387_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0851_),
    .B1(_0876_),
    .B2(\u_cpu.cpu.immdec.imm24_20[3] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1388_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_0875_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1389_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0851_),
    .B1(_0876_),
    .B2(\u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1390_ (.A1(_0877_),
    .A2(_0878_),
    .A3(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1391_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_0874_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1392_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_0859_),
    .A4(_0866_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1393_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_0862_),
    .A3(_0881_),
    .A4(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1394_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .B(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1395_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0851_),
    .B1(_0876_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1396_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A3(_0871_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1397_ (.A1(_0865_),
    .A2(_0868_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1398_ (.A1(_0886_),
    .A2(_0887_),
    .B(_0851_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1399_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_0851_),
    .B1(_0876_),
    .B2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .C(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1400_ (.A1(_0884_),
    .A2(_0885_),
    .A3(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1401_ (.A1(_0880_),
    .A2(_0890_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1402_ (.I(_0851_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1403_ (.I(io_in[1]),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1404_ (.I(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1405_ (.A1(_0892_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1406_ (.I(_0893_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1407_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1408_ (.I(_0895_),
    .Z(\u_arbiter.o_wb_cpu_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1409_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0894_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1410_ (.I(_0896_),
    .Z(\u_arbiter.o_wb_cpu_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1411_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1412_ (.I(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1413_ (.I(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1414_ (.I(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1415_ (.A1(_0900_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1416_ (.A1(_0900_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1417_ (.A1(_0894_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1418_ (.A1(_0892_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1419_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1420_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1421_ (.A1(_0901_),
    .A2(_0903_),
    .B(_0906_),
    .ZN(\u_arbiter.o_wb_cpu_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1422_ (.I(_0904_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1423_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0902_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1424_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .A2(_0905_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1425_ (.A1(_0907_),
    .A2(_0908_),
    .B(_0909_),
    .ZN(\u_arbiter.o_wb_cpu_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1426_ (.A1(_0900_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1427_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1428_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .A2(_0905_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1429_ (.A1(_0907_),
    .A2(_0911_),
    .B(_0912_),
    .ZN(\u_arbiter.o_wb_cpu_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1430_ (.A1(_0897_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1431_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1432_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .A2(_0905_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1433_ (.A1(_0907_),
    .A2(_0914_),
    .B(_0915_),
    .ZN(\u_arbiter.o_wb_cpu_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1434_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_0913_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1435_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A3(_0913_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1436_ (.A1(_0894_),
    .A2(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1437_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .A2(_0905_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1438_ (.A1(_0916_),
    .A2(_0918_),
    .B(_0919_),
    .ZN(\u_arbiter.o_wb_cpu_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1439_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0917_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1440_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .A2(_0905_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1441_ (.A1(_0907_),
    .A2(_0920_),
    .B(_0921_),
    .ZN(\u_arbiter.o_wb_cpu_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1442_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1443_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_0913_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1444_ (.A1(_0922_),
    .A2(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1445_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1446_ (.I(_0904_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1447_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1448_ (.A1(_0905_),
    .A2(_0924_),
    .A3(_0925_),
    .B(_0927_),
    .ZN(\u_arbiter.o_wb_cpu_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1449_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0925_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1450_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1451_ (.A1(_0929_),
    .A2(_0922_),
    .A3(_0923_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1452_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .A2(_0926_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1453_ (.A1(_0905_),
    .A2(_0928_),
    .A3(_0930_),
    .B(_0931_),
    .ZN(\u_arbiter.o_wb_cpu_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1454_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .A2(_0905_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1455_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0930_),
    .B(_0904_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1456_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0930_),
    .B(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1457_ (.A1(_0932_),
    .A2(_0934_),
    .ZN(\u_arbiter.o_wb_cpu_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1458_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0930_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1459_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1460_ (.A1(_0929_),
    .A2(_0922_),
    .A3(_0923_),
    .A4(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1461_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .A2(_0926_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1462_ (.A1(_0905_),
    .A2(_0935_),
    .A3(_0937_),
    .B(_0938_),
    .ZN(\u_arbiter.o_wb_cpu_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1463_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_0937_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1464_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_0905_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1465_ (.A1(_0907_),
    .A2(_0939_),
    .B(_0940_),
    .ZN(\u_arbiter.o_wb_cpu_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1466_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_0937_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1467_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_0937_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1468_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_0926_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1469_ (.A1(_0905_),
    .A2(_0941_),
    .A3(_0942_),
    .B(_0943_),
    .ZN(\u_arbiter.o_wb_cpu_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1470_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .A2(_0905_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1471_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0942_),
    .B(_0904_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1472_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0942_),
    .B(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1473_ (.A1(_0944_),
    .A2(_0946_),
    .ZN(\u_arbiter.o_wb_cpu_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1474_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0942_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1475_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1476_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_0937_),
    .A4(_0948_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1477_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .A2(_0926_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1478_ (.A1(_0905_),
    .A2(_0947_),
    .A3(_0949_),
    .B(_0950_),
    .ZN(\u_arbiter.o_wb_cpu_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1479_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0949_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1480_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(_0951_),
    .S(_0894_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1481_ (.I(_0952_),
    .Z(\u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1482_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0949_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1483_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A3(_0949_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1484_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_0904_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1485_ (.A1(_0905_),
    .A2(_0953_),
    .A3(_0954_),
    .B(_0955_),
    .ZN(\u_arbiter.o_wb_cpu_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1486_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0954_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1487_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(_0956_),
    .S(_0894_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1488_ (.I(_0957_),
    .Z(\u_arbiter.o_wb_cpu_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1489_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1490_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A4(_0949_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1491_ (.A1(_0958_),
    .A2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1492_ (.A1(_0958_),
    .A2(_0959_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1493_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_0904_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1494_ (.A1(_0905_),
    .A2(_0960_),
    .A3(_0961_),
    .B(_0962_),
    .ZN(\u_arbiter.o_wb_cpu_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1495_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0960_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1496_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .A2(_0926_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1497_ (.A1(_0907_),
    .A2(_0963_),
    .B(_0964_),
    .ZN(\u_arbiter.o_wb_cpu_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1498_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0960_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1499_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1500_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .A2(_0926_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1501_ (.A1(_0907_),
    .A2(_0966_),
    .B(_0967_),
    .ZN(\u_arbiter.o_wb_cpu_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1502_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A3(_0960_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1503_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1504_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .A2(_0926_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1505_ (.A1(_0907_),
    .A2(_0969_),
    .B(_0970_),
    .ZN(\u_arbiter.o_wb_cpu_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1506_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A4(_0960_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1507_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1508_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_0926_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1509_ (.A1(_0907_),
    .A2(_0972_),
    .B(_0973_),
    .ZN(\u_arbiter.o_wb_cpu_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1510_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0971_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1511_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1512_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_0926_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1513_ (.A1(_0907_),
    .A2(_0975_),
    .B(_0976_),
    .ZN(\u_arbiter.o_wb_cpu_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1514_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A3(_0971_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1515_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0977_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1516_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_0926_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1517_ (.A1(_0907_),
    .A2(_0978_),
    .B(_0979_),
    .ZN(\u_arbiter.o_wb_cpu_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1518_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A4(_0971_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1519_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1520_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .A2(_0926_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1521_ (.A1(_0907_),
    .A2(_0981_),
    .B(_0982_),
    .ZN(\u_arbiter.o_wb_cpu_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1522_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0980_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1523_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_0983_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1524_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_0926_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1525_ (.A1(_0907_),
    .A2(_0984_),
    .B(_0985_),
    .ZN(\u_arbiter.o_wb_cpu_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1526_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A3(_0980_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1527_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1528_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_0926_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1529_ (.A1(_0907_),
    .A2(_0987_),
    .B(_0988_),
    .ZN(\u_arbiter.o_wb_cpu_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1530_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A4(_0980_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1531_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1532_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_0926_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1533_ (.A1(_0907_),
    .A2(_0990_),
    .B(_0991_),
    .ZN(\u_arbiter.o_wb_cpu_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1534_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0989_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1535_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A3(_0989_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1536_ (.A1(_0894_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1537_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_0926_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1538_ (.A1(_0992_),
    .A2(_0994_),
    .B(_0995_),
    .ZN(\u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1539_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0993_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1540_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A2(_0894_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1541_ (.A1(_0894_),
    .A2(_0996_),
    .B(_0997_),
    .ZN(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1542_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1543_ (.A1(\u_cpu.rf_ram_if.wen1_r ),
    .A2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1544_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0849_),
    .A3(_0850_),
    .A4(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1545_ (.A1(_0999_),
    .A2(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1546_ (.I(_1001_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1547_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1548_ (.A1(_0858_),
    .A2(_0861_),
    .A3(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1549_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1550_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1551_ (.A1(\u_cpu.rf_ram.data[0] ),
    .A2(_0999_),
    .A3(_1000_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1552_ (.I(_0999_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1553_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0849_),
    .A3(_0850_),
    .A4(\u_cpu.rf_ram_if.wen0_r ),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1554_ (.A1(_1007_),
    .A2(_1008_),
    .B(\u_cpu.rf_ram.rdata[0] ),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1555_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1556_ (.I(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1557_ (.A1(_1006_),
    .A2(_1009_),
    .B(\u_cpu.rf_ram.regzero ),
    .C(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1558_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(_1011_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1559_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1560_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1561_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1562_ (.A1(_0855_),
    .A2(_1016_),
    .A3(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1563_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1015_),
    .A3(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1564_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1017_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1565_ (.A1(_0855_),
    .A2(\u_cpu.cpu.branch_op ),
    .A3(_0853_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1566_ (.A1(_1014_),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1567_ (.A1(_1014_),
    .A2(_1018_),
    .A3(_1019_),
    .B(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1568_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1569_ (.A1(_1005_),
    .A2(_1012_),
    .A3(_1013_),
    .B(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1570_ (.A1(_1003_),
    .A2(_1024_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1571_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1572_ (.A1(_1004_),
    .A2(_1025_),
    .B(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1573_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1574_ (.I(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1575_ (.I0(_1003_),
    .I1(_1027_),
    .S(_1029_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1576_ (.I(_1030_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1577_ (.I(_0860_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1578_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1579_ (.A1(_0853_),
    .A2(\u_cpu.cpu.csr_imm ),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1580_ (.A1(_0853_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1581_ (.A1(_1031_),
    .A2(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1582_ (.A1(_1012_),
    .A2(_1013_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1583_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1584_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1585_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_0867_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1586_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_1037_),
    .A3(_1038_),
    .A4(_1039_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1587_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1588_ (.A1(_1014_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1589_ (.A1(_1041_),
    .A2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1590_ (.A1(_0864_),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_0867_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1591_ (.A1(_1029_),
    .A2(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1592_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .A2(_1041_),
    .B(_1043_),
    .C(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1593_ (.I(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1594_ (.A1(_0868_),
    .A2(_1036_),
    .B1(_1040_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1595_ (.A1(_0860_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .B(_1034_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1596_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_1035_),
    .B1(_1048_),
    .B2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1597_ (.A1(_0886_),
    .A2(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1598_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_0873_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1599_ (.A1(_1051_),
    .A2(_1052_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1600_ (.I(_0852_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1601_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.init_done ),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1602_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A3(_0857_),
    .A4(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1603_ (.A1(_0860_),
    .A2(_0853_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1604_ (.A1(\u_cpu.cpu.branch_op ),
    .A2(_1016_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1605_ (.A1(_0861_),
    .A2(_1056_),
    .A3(_1057_),
    .B(_0855_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1606_ (.A1(_1029_),
    .A2(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1607_ (.A1(_1055_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1608_ (.A1(_0860_),
    .A2(_0856_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1609_ (.A1(_0853_),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .B(_1061_),
    .C(\u_cpu.cpu.state.init_done ),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1610_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1611_ (.A1(_1060_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1612_ (.A1(_1053_),
    .A2(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1613_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_1038_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1614_ (.A1(_0857_),
    .A2(\u_arbiter.i_wb_cpu_dbus_we ),
    .B1(_0863_),
    .B2(_0870_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1615_ (.A1(_1016_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1616_ (.A1(_1017_),
    .A2(_1067_),
    .A3(_1068_),
    .B(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1617_ (.I(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1618_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1619_ (.A1(_1055_),
    .A2(_1059_),
    .B1(_1062_),
    .B2(\u_cpu.cpu.state.stage_two_req ),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1620_ (.I(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1621_ (.A1(_0852_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1622_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1623_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_1075_),
    .B(_1022_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1624_ (.A1(_0855_),
    .A2(_1016_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1625_ (.A1(_0857_),
    .A2(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1626_ (.I0(_1074_),
    .I1(_1076_),
    .S(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1627_ (.A1(_1071_),
    .A2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1628_ (.A1(_1066_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1629_ (.A1(_0857_),
    .A2(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1630_ (.A1(_0857_),
    .A2(_1065_),
    .B(_1082_),
    .C(_0873_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1631_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1632_ (.A1(_1084_),
    .A2(_1003_),
    .A3(_1024_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1633_ (.A1(_0866_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1634_ (.A1(_0860_),
    .A2(_1032_),
    .A3(_1024_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1635_ (.A1(_1032_),
    .A2(_1024_),
    .B(\u_cpu.cpu.bne_or_bge ),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1636_ (.A1(_1032_),
    .A2(_1024_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1637_ (.A1(_0853_),
    .A2(_1087_),
    .A3(_1088_),
    .A4(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1638_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_1038_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1639_ (.A1(_0860_),
    .A2(_0854_),
    .A3(\u_cpu.cpu.alu.cmp_r ),
    .A4(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1640_ (.A1(_1074_),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1641_ (.A1(_0856_),
    .A2(_1057_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1642_ (.A1(_1086_),
    .A2(_1090_),
    .A3(_1093_),
    .B(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1643_ (.A1(_1078_),
    .A2(_1066_),
    .A3(_1080_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1644_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1645_ (.A1(_1031_),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B1(\u_cpu.cpu.mem_bytecnt[0] ),
    .B2(_0861_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1646_ (.I0(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(_0852_),
    .S1(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1647_ (.A1(_1098_),
    .A2(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1648_ (.A1(_1097_),
    .A2(_1098_),
    .B(_1100_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1649_ (.A1(_0853_),
    .A2(_1100_),
    .B(_0855_),
    .C(_1016_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1650_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1651_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1652_ (.A1(_1102_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_1041_),
    .C(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1653_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1654_ (.A1(_1104_),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1655_ (.A1(_0857_),
    .A2(_1016_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1656_ (.A1(_1106_),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1657_ (.A1(_0041_),
    .A2(_1101_),
    .B(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1658_ (.A1(_1048_),
    .A2(_1095_),
    .A3(_1096_),
    .A4(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1659_ (.A1(_0886_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1660_ (.A1(_1083_),
    .A2(_1111_),
    .ZN(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1661_ (.A1(_1006_),
    .A2(_1009_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1662_ (.I0(\u_cpu.rf_ram.rdata[1] ),
    .I1(\u_cpu.rf_ram.data[1] ),
    .S(_0026_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1663_ (.I(_1112_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1664_ (.I0(\u_cpu.rf_ram.rdata[2] ),
    .I1(\u_cpu.rf_ram.data[2] ),
    .S(_0026_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1665_ (.I(_1113_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1666_ (.I0(\u_cpu.rf_ram.rdata[3] ),
    .I1(\u_cpu.rf_ram.data[3] ),
    .S(_0026_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1667_ (.I(_1114_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1668_ (.I0(\u_cpu.rf_ram.rdata[4] ),
    .I1(\u_cpu.rf_ram.data[4] ),
    .S(_0026_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1669_ (.I(_1115_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1670_ (.I0(\u_cpu.rf_ram.rdata[5] ),
    .I1(\u_cpu.rf_ram.data[5] ),
    .S(_0026_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1671_ (.I(_1116_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1672_ (.I0(\u_cpu.rf_ram.rdata[6] ),
    .I1(\u_cpu.rf_ram.data[6] ),
    .S(_0026_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1673_ (.I(_1117_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1674_ (.I0(\u_cpu.rf_ram.rdata[7] ),
    .I1(\u_cpu.rf_ram.data[7] ),
    .S(_0026_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1675_ (.I(_1118_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1676_ (.I0(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .S(_0998_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1677_ (.I(_1119_),
    .Z(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1678_ (.I0(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .S(_0998_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1679_ (.I(_1120_),
    .Z(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1680_ (.I0(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .S(_0998_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1681_ (.I(_1121_),
    .Z(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1682_ (.I0(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .S(_0998_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1683_ (.I(_1122_),
    .Z(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1684_ (.I0(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .S(_0998_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1685_ (.I(_1123_),
    .Z(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1686_ (.I0(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .S(_0998_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1687_ (.I(_1124_),
    .Z(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1688_ (.I0(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .S(_0998_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1689_ (.I(_1125_),
    .Z(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1690_ (.I(_0998_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1691_ (.I0(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .I1(\u_cpu.cpu.o_wdata0 ),
    .S(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1692_ (.I(_1127_),
    .Z(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1693_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1694_ (.A1(_1128_),
    .A2(_0018_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1695_ (.I0(\u_cpu.rf_ram_if.rdata1[1] ),
    .I1(_1129_),
    .S(_1010_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1696_ (.I(_1130_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1697_ (.A1(_1128_),
    .A2(_0019_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1698_ (.I0(\u_cpu.rf_ram_if.rdata1[2] ),
    .I1(_1131_),
    .S(_1010_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1699_ (.I(_1132_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1700_ (.A1(_1128_),
    .A2(_0020_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1701_ (.I0(\u_cpu.rf_ram_if.rdata1[3] ),
    .I1(_1133_),
    .S(_1010_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1702_ (.I(_1134_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1703_ (.A1(_1128_),
    .A2(_0021_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1704_ (.I0(\u_cpu.rf_ram_if.rdata1[4] ),
    .I1(_1135_),
    .S(_1010_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1705_ (.I(_1136_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1706_ (.A1(_1128_),
    .A2(_0022_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1707_ (.I0(\u_cpu.rf_ram_if.rdata1[5] ),
    .I1(_1137_),
    .S(_1010_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1708_ (.I(_1138_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1709_ (.A1(_1128_),
    .A2(_0023_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1710_ (.I0(\u_cpu.rf_ram_if.rdata1[6] ),
    .I1(_1139_),
    .S(_1010_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1711_ (.I(_1140_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1712_ (.A1(_1006_),
    .A2(_1009_),
    .B(\u_cpu.rf_ram.regzero ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1713_ (.I0(\u_cpu.rf_ram_if.rdata0[1] ),
    .I1(_1141_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1714_ (.I(_1142_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1715_ (.I0(\u_cpu.rf_ram_if.rdata0[2] ),
    .I1(_1129_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1716_ (.I(_1143_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1717_ (.I0(\u_cpu.rf_ram_if.rdata0[3] ),
    .I1(_1131_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1718_ (.I(_1144_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1719_ (.I0(\u_cpu.rf_ram_if.rdata0[4] ),
    .I1(_1133_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1720_ (.I(_1145_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1721_ (.I0(\u_cpu.rf_ram_if.rdata0[5] ),
    .I1(_1135_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1722_ (.I(_1146_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1723_ (.I0(\u_cpu.rf_ram_if.rdata0[6] ),
    .I1(_1137_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1724_ (.I(_1147_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1725_ (.I0(\u_cpu.rf_ram_if.rdata0[7] ),
    .I1(_1139_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1726_ (.I(_1148_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1727_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1728_ (.A1(_1001_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1729_ (.A1(\u_cpu.raddr[0] ),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1730_ (.I(_1151_),
    .Z(\u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1731_ (.A1(\u_cpu.raddr[0] ),
    .A2(_1150_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1732_ (.A1(\u_cpu.raddr[1] ),
    .A2(_1152_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1733_ (.I(_1153_),
    .Z(\u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1734_ (.A1(_0865_),
    .A2(_0886_),
    .B(_1126_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1735_ (.A1(\u_cpu.cpu.immdec.imm11_7[0] ),
    .A2(_0998_),
    .A3(_0873_),
    .B(_1001_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1736_ (.A1(_0889_),
    .A2(_1001_),
    .B1(_1154_),
    .B2(_1155_),
    .ZN(\u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1737_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_0998_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1738_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_1126_),
    .B(_0026_),
    .C(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1739_ (.A1(_0884_),
    .A2(_0026_),
    .B1(_1157_),
    .B2(_0886_),
    .ZN(\u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1740_ (.A1(_1126_),
    .A2(_0886_),
    .A3(_1001_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1741_ (.I(\u_cpu.cpu.immdec.imm11_7[2] ),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1742_ (.A1(_0885_),
    .A2(_1001_),
    .B1(_1158_),
    .B2(_1159_),
    .ZN(\u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1743_ (.I(_1158_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1744_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1745_ (.A1(_0877_),
    .A2(_1001_),
    .B(_1161_),
    .ZN(\u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1746_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1747_ (.A1(_0879_),
    .A2(_1001_),
    .B1(_1158_),
    .B2(_1162_),
    .ZN(\u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1748_ (.A1(_0878_),
    .A2(_0026_),
    .B(_1160_),
    .ZN(\u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1749_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1750_ (.A1(_1031_),
    .A2(_1163_),
    .B1(_0861_),
    .B2(_1053_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1751_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1752_ (.A1(_0855_),
    .A2(_0857_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1753_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_1165_),
    .A3(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1754_ (.A1(_1164_),
    .A2(_1167_),
    .B(_0907_),
    .ZN(\u_arbiter.o_wb_cpu_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1755_ (.A1(_1005_),
    .A2(_0894_),
    .ZN(\u_arbiter.o_wb_cpu_we ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1756_ (.A1(_0857_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1757_ (.I(_1016_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1758_ (.A1(_0857_),
    .A2(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1759_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.bufreg.c_r ),
    .A3(_1168_),
    .A4(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1760_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_1168_),
    .A3(_1170_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1761_ (.A1(\u_cpu.cpu.bufreg.c_r ),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1762_ (.A1(_1016_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1763_ (.A1(_1174_),
    .A2(_1068_),
    .B(_1091_),
    .C(_0857_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1764_ (.A1(_0856_),
    .A2(_1022_),
    .A3(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1765_ (.A1(_1173_),
    .A2(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1766_ (.A1(_1171_),
    .A2(_1177_),
    .B(_1064_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1767_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1070_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1768_ (.A1(_1078_),
    .A2(_1076_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1769_ (.A1(_1078_),
    .A2(_1065_),
    .B(_1179_),
    .C(_1071_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1770_ (.A1(_1054_),
    .A2(_1058_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1771_ (.A1(_1029_),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1772_ (.A1(_1178_),
    .A2(_1180_),
    .B(_1182_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1773_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1774_ (.A1(_1104_),
    .A2(_1105_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1775_ (.A1(_1183_),
    .A2(_1184_),
    .B(_1182_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1776_ (.A1(_0874_),
    .A2(_1165_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1777_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A3(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1778_ (.A1(_1016_),
    .A2(\u_arbiter.i_wb_cpu_dbus_we ),
    .B(_1107_),
    .C(_0856_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1779_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_1185_),
    .B(_1186_),
    .C(_1181_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1780_ (.A1(_0886_),
    .A2(_1187_),
    .B(_1165_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1781_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_0852_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1782_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_1188_),
    .B(_1031_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1783_ (.A1(_0852_),
    .A2(_1163_),
    .B(_1031_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1784_ (.A1(_1163_),
    .A2(_1188_),
    .B(_1031_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1785_ (.I(_0897_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1786_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_0894_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1787_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1788_ (.I(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1789_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1790_ (.A1(_0891_),
    .A2(_1193_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(_1031_),
    .A2(_0855_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1792_ (.A1(_1054_),
    .A2(_1058_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1793_ (.A1(_1194_),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1794_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A4(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1795_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1796_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1797_ (.A1(_1014_),
    .A2(_1061_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1798_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_1200_),
    .B(_1196_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1799_ (.A1(_1196_),
    .A2(_1199_),
    .B(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1800_ (.A1(_0860_),
    .A2(_0854_),
    .A3(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1801_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_0904_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1802_ (.A1(_0856_),
    .A2(_1203_),
    .B(_1204_),
    .C(_0858_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1803_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_0869_),
    .A3(_1165_),
    .A4(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1804_ (.A1(_1193_),
    .A2(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1805_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_1207_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1806_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1807_ (.A1(_0215_),
    .A2(_0849_),
    .A3(_0850_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1808_ (.A1(_1149_),
    .A2(_1207_),
    .A3(_0216_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1809_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1810_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0216_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1811_ (.A1(_1193_),
    .A2(_1206_),
    .A3(_0217_),
    .A4(_0218_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1812_ (.I(_0219_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1813_ (.A1(\u_cpu.raddr[1] ),
    .A2(_0217_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1814_ (.A1(_1207_),
    .A2(_0220_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1815_ (.A1(_1014_),
    .A2(_1195_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1816_ (.A1(_0891_),
    .A2(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1817_ (.I(_0222_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1818_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1819_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1820_ (.A1(_0891_),
    .A2(_0223_),
    .A3(_0224_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1821_ (.A1(\u_cpu.cpu.mem_bytecnt[0] ),
    .A2(_0224_),
    .B(_0892_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1822_ (.A1(\u_cpu.cpu.mem_bytecnt[0] ),
    .A2(_0224_),
    .B(_0225_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1823_ (.A1(\u_cpu.cpu.mem_bytecnt[0] ),
    .A2(_0224_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1824_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1825_ (.A1(_0891_),
    .A2(_0227_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1826_ (.A1(_0891_),
    .A2(_1014_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1827_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_0228_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1828_ (.I(\u_cpu.rf_ram_if.rgnt ),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1829_ (.A1(_0230_),
    .A2(_1206_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1830_ (.A1(_0892_),
    .A2(_1165_),
    .A3(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1831_ (.A1(_0229_),
    .A2(_0232_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1832_ (.A1(_0892_),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1833_ (.I(_0233_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1834_ (.A1(_0891_),
    .A2(_1102_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1835_ (.A1(_0892_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1836_ (.I(_0234_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1837_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_0228_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1838_ (.A1(_1164_),
    .A2(_1166_),
    .A3(_0032_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1839_ (.A1(_0235_),
    .A2(_0236_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1840_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_0228_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1841_ (.A1(_0860_),
    .A2(_0853_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1842_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_0853_),
    .B(_0860_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1843_ (.A1(_1032_),
    .A2(_1024_),
    .B(_0239_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1844_ (.A1(_1032_),
    .A2(_1024_),
    .B(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1845_ (.A1(_1027_),
    .A2(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1846_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_1091_),
    .B(_1085_),
    .C(_0238_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1847_ (.A1(_0238_),
    .A2(_0242_),
    .B(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1848_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_0244_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1849_ (.A1(_1016_),
    .A2(_0245_),
    .B(_0032_),
    .C(_0857_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1850_ (.A1(_0237_),
    .A2(_0246_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1851_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_1075_),
    .A3(_0039_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1852_ (.I(_0247_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1853_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_0228_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1854_ (.A1(_0891_),
    .A2(_0221_),
    .B(_0248_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1855_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B(\u_cpu.cpu.mem_bytecnt[0] ),
    .C(_0852_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1856_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1857_ (.A1(_1029_),
    .A2(_0249_),
    .A3(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1858_ (.A1(_1194_),
    .A2(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1859_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(_1196_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1860_ (.A1(_0252_),
    .A2(_0253_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1861_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(_1196_),
    .B(_1204_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1862_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_0904_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1863_ (.I(_0256_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1864_ (.A1(_0257_),
    .A2(_0252_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1865_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1866_ (.A1(_0254_),
    .A2(_0255_),
    .B(_0259_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1867_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_1196_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1868_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .B(_1196_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1869_ (.A1(_0252_),
    .A2(_0261_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1870_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(_0254_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1871_ (.A1(_0260_),
    .A2(_0262_),
    .B(_1204_),
    .C(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1872_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_1204_),
    .B(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1873_ (.I(_0265_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1874_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_1196_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1875_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .B(_1196_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1876_ (.A1(_0252_),
    .A2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1877_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_0262_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1878_ (.A1(_0266_),
    .A2(_0268_),
    .B(_1204_),
    .C(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1879_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_1204_),
    .B(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1880_ (.I(_0271_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1881_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1882_ (.I(_0257_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1883_ (.A1(_1196_),
    .A2(_1197_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1884_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_1196_),
    .B(_0252_),
    .C(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1885_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_0268_),
    .B(_0257_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1886_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0275_),
    .B2(_0276_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1887_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_1197_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1888_ (.A1(_1196_),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1889_ (.A1(_1204_),
    .A2(_0252_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1890_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1891_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_1196_),
    .B1(_1198_),
    .B2(_0278_),
    .C(_0280_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1892_ (.I(_0258_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1893_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1894_ (.A1(_0281_),
    .A2(_0283_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1895_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_0273_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1896_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0258_),
    .B1(_0280_),
    .B2(_1202_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1897_ (.A1(_0284_),
    .A2(_0285_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1898_ (.I(_0280_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1899_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .A2(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1900_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1901_ (.A1(_0287_),
    .A2(_0288_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1902_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1903_ (.I(_0289_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1904_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_0286_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1905_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1906_ (.A1(_0290_),
    .A2(_0291_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1907_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1908_ (.I(_0292_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_0286_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1910_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1911_ (.A1(_0293_),
    .A2(_0294_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1912_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_0286_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1913_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1914_ (.A1(_0295_),
    .A2(_0296_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1915_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1916_ (.I(_0297_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1917_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_0286_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1918_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1919_ (.A1(_0298_),
    .A2(_0299_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1920_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .A2(_0286_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1921_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1922_ (.A1(_0300_),
    .A2(_0301_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1923_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_0286_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1924_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1925_ (.A1(_0302_),
    .A2(_0303_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1926_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1927_ (.I(_0304_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1928_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(_0286_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1929_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1930_ (.A1(_0305_),
    .A2(_0306_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1931_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_0286_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1932_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1933_ (.A1(_0307_),
    .A2(_0308_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1934_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_0286_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1935_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_0273_),
    .B1(_0282_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1936_ (.A1(_0309_),
    .A2(_0310_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1937_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_0286_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1938_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_0273_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1939_ (.A1(_0311_),
    .A2(_0312_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1940_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .A2(_0286_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1941_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_0273_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1942_ (.A1(_0313_),
    .A2(_0314_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1943_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1944_ (.I(_0315_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1945_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0280_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1946_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_0273_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1947_ (.A1(_0316_),
    .A2(_0317_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1948_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0282_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1949_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_0257_),
    .B1(_0280_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1950_ (.A1(_0318_),
    .A2(_0319_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1951_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1952_ (.I(_0320_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1953_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1954_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1955_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_1204_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1956_ (.A1(_0321_),
    .A2(_0282_),
    .B1(_0286_),
    .B2(_0322_),
    .C(_0323_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1957_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1958_ (.I(_0324_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1959_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .C1(_0280_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1960_ (.I(_0325_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1961_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1962_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1963_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_1204_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1964_ (.A1(_0326_),
    .A2(_0282_),
    .B1(_0286_),
    .B2(_0327_),
    .C(_0328_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1965_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1966_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_1204_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1967_ (.A1(_0327_),
    .A2(_0282_),
    .B1(_0286_),
    .B2(_0329_),
    .C(_0330_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1968_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_1204_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1969_ (.A1(_0329_),
    .A2(_0282_),
    .B1(_0286_),
    .B2(_1024_),
    .C(_0331_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1970_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1971_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_0894_),
    .A3(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1972_ (.I(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1973_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0897_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1974_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0897_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1975_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0897_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1976_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0897_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1977_ (.A1(_0335_),
    .A2(_0336_),
    .A3(_0337_),
    .A4(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1978_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_0899_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1979_ (.A1(_0339_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1980_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0898_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1981_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1982_ (.A1(_0341_),
    .A2(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1983_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0899_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1984_ (.A1(_0899_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1985_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1986_ (.A1(_0345_),
    .A2(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1987_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1988_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[6] ),
    .B(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1989_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1990_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1991_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1992_ (.A1(_0899_),
    .A2(_0272_),
    .B(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1993_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0898_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1994_ (.I0(\u_arbiter.i_wb_cpu_rdt[2] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0898_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1995_ (.A1(_0354_),
    .A2(_0355_),
    .A3(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1996_ (.A1(_0350_),
    .A2(_0352_),
    .A3(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1997_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1998_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1999_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_0898_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2000_ (.A1(_0360_),
    .A2(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2001_ (.A1(_0358_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2002_ (.A1(_0348_),
    .A2(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2003_ (.A1(_0344_),
    .A2(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2004_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2005_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2006_ (.I0(\u_arbiter.i_wb_cpu_rdt[1] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_0899_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2007_ (.A1(_0367_),
    .A2(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2008_ (.A1(_0360_),
    .A2(_0361_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2009_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_0898_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2010_ (.A1(_0370_),
    .A2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2011_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2012_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2013_ (.A1(_0339_),
    .A2(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2014_ (.A1(_0372_),
    .A2(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2015_ (.A1(_0360_),
    .A2(_0371_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2016_ (.A1(_0376_),
    .A2(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2017_ (.A1(_0367_),
    .A2(_0347_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2018_ (.A1(_0345_),
    .A2(_0368_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2019_ (.A1(_0362_),
    .A2(_0379_),
    .B(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2020_ (.I(_0333_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2021_ (.A1(_0369_),
    .A2(_0378_),
    .B1(_0381_),
    .B2(_0356_),
    .C(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2022_ (.A1(_1169_),
    .A2(_0334_),
    .B1(_0365_),
    .B2(_0383_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2023_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0898_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2024_ (.I(_0384_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2025_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2026_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2027_ (.A1(_0385_),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2028_ (.A1(_0369_),
    .A2(_0388_),
    .B1(_0381_),
    .B2(_0354_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2029_ (.A1(\u_cpu.cpu.decode.opcode[1] ),
    .A2(_0334_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2030_ (.A1(_0334_),
    .A2(_0389_),
    .B(_0390_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2031_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2032_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2033_ (.A1(_0360_),
    .A2(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2034_ (.A1(_0388_),
    .A2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2035_ (.A1(_0333_),
    .A2(_0381_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2036_ (.A1(_0367_),
    .A2(_0394_),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2037_ (.I(_0392_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2038_ (.A1(_0397_),
    .A2(_0358_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2039_ (.A1(_0367_),
    .A2(_0385_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2040_ (.A1(_0344_),
    .A2(_0347_),
    .A3(_0398_),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2041_ (.A1(_0385_),
    .A2(_0397_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2042_ (.A1(_0345_),
    .A2(_0368_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2043_ (.A1(_0367_),
    .A2(_0347_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2044_ (.A1(_0401_),
    .A2(_0402_),
    .B(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2045_ (.A1(_0333_),
    .A2(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2046_ (.A1(_0855_),
    .A2(_0334_),
    .B1(_0355_),
    .B2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2047_ (.A1(_0396_),
    .A2(_0400_),
    .B(_0406_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2048_ (.I(_1192_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2049_ (.A1(_0345_),
    .A2(_0347_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2050_ (.A1(_0362_),
    .A2(_0371_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2051_ (.A1(_0899_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2052_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[11] ),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2053_ (.A1(_0898_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2054_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[10] ),
    .B(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2055_ (.A1(_0411_),
    .A2(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2056_ (.A1(_0409_),
    .A2(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2057_ (.A1(_0376_),
    .A2(_0394_),
    .A3(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2058_ (.A1(_0367_),
    .A2(_0397_),
    .B1(_0352_),
    .B2(_0381_),
    .C(_0382_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2059_ (.A1(_0408_),
    .A2(_0416_),
    .B(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2060_ (.A1(_1005_),
    .A2(_0407_),
    .B(_0418_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2061_ (.A1(_0385_),
    .A2(_0361_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2062_ (.A1(_0377_),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2063_ (.A1(_1192_),
    .A2(_0404_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2064_ (.A1(_0345_),
    .A2(_0420_),
    .B(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2065_ (.A1(_0857_),
    .A2(_1192_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2066_ (.A1(_0364_),
    .A2(_0422_),
    .B1(_0405_),
    .B2(_0350_),
    .C(_0423_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2067_ (.I(\u_cpu.cpu.bne_or_bge ),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2068_ (.A1(_0372_),
    .A2(_0375_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2069_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_0899_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2070_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_0899_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2071_ (.A1(_0426_),
    .A2(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2072_ (.A1(_0401_),
    .A2(_0387_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2073_ (.A1(_0414_),
    .A2(_0428_),
    .B(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2074_ (.A1(_0356_),
    .A2(_0425_),
    .B1(_0393_),
    .B2(_0371_),
    .C(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2075_ (.A1(_0408_),
    .A2(_0377_),
    .B(_0404_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2076_ (.A1(_0385_),
    .A2(_0361_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2077_ (.A1(_0343_),
    .A2(_0432_),
    .B1(_0433_),
    .B2(_0348_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2078_ (.A1(_0408_),
    .A2(_0431_),
    .B(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2079_ (.A1(_0407_),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2080_ (.A1(_0424_),
    .A2(_0407_),
    .B(_0436_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2081_ (.A1(_0336_),
    .A2(_0350_),
    .B(_0411_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2082_ (.A1(_0343_),
    .A2(_0388_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2083_ (.A1(_0354_),
    .A2(_0425_),
    .B1(_0409_),
    .B2(_0437_),
    .C(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2084_ (.A1(_0408_),
    .A2(_0439_),
    .B(_0399_),
    .C(_0404_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2085_ (.A1(_0371_),
    .A2(_0404_),
    .B(_0440_),
    .C(_1192_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2086_ (.A1(_1031_),
    .A2(_0407_),
    .B(_0441_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2087_ (.A1(_0350_),
    .A2(_0352_),
    .A3(_0414_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2088_ (.A1(_0355_),
    .A2(_0425_),
    .B1(_0409_),
    .B2(_0442_),
    .C(_0438_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2089_ (.A1(_0360_),
    .A2(_0380_),
    .B1(_0443_),
    .B2(_0408_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2090_ (.A1(_0407_),
    .A2(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2091_ (.A1(_0854_),
    .A2(_0407_),
    .B(_0445_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2092_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_0900_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2093_ (.A1(_0356_),
    .A2(_0387_),
    .A3(_0419_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2094_ (.A1(_0343_),
    .A2(_0425_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2095_ (.A1(_0438_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2096_ (.A1(_0345_),
    .A2(_0447_),
    .A3(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2097_ (.A1(_0385_),
    .A2(_0397_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2098_ (.A1(_0344_),
    .A2(_0363_),
    .B1(_0451_),
    .B2(_0356_),
    .C(_0347_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2099_ (.A1(_0356_),
    .A2(_0393_),
    .B(_0379_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2100_ (.A1(_0333_),
    .A2(_0403_),
    .A3(_0452_),
    .A4(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2101_ (.A1(_0405_),
    .A2(_0446_),
    .B1(_0450_),
    .B2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2102_ (.A1(_0863_),
    .A2(_0407_),
    .B(_0455_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2103_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_0900_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2104_ (.A1(_0397_),
    .A2(_0387_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2105_ (.A1(_0385_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2106_ (.A1(_0354_),
    .A2(_0458_),
    .B(_0448_),
    .C(_0367_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2107_ (.A1(_0367_),
    .A2(_0354_),
    .A3(_0451_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2108_ (.A1(_0368_),
    .A2(_0459_),
    .B(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(_0354_),
    .A2(_0393_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2110_ (.A1(_0402_),
    .A2(_0462_),
    .B(_0421_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2111_ (.A1(_0405_),
    .A2(_0456_),
    .B1(_0461_),
    .B2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2112_ (.A1(_0864_),
    .A2(_0407_),
    .B(_0464_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2113_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_0899_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2114_ (.A1(_0899_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2115_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[4] ),
    .B(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2116_ (.A1(_0369_),
    .A2(_0448_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2117_ (.A1(_0448_),
    .A2(_0458_),
    .B(_0369_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2118_ (.A1(_0367_),
    .A2(_0368_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2119_ (.A1(_0467_),
    .A2(_0468_),
    .B1(_0469_),
    .B2(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2120_ (.I(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2121_ (.A1(_0355_),
    .A2(_0393_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2122_ (.A1(_0397_),
    .A2(_0426_),
    .B1(_0401_),
    .B2(_0465_),
    .C(_0379_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2123_ (.A1(_0379_),
    .A2(_0472_),
    .B1(_0473_),
    .B2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2124_ (.A1(_0405_),
    .A2(_0465_),
    .B1(_0475_),
    .B2(_0395_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2125_ (.A1(_1037_),
    .A2(_0407_),
    .B(_0476_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2126_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_0334_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2127_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_0899_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2128_ (.A1(_0387_),
    .A2(_0433_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2129_ (.A1(_0343_),
    .A2(_0479_),
    .B(_0369_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2130_ (.A1(_0343_),
    .A2(_0385_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2131_ (.A1(_0335_),
    .A2(_0413_),
    .A3(_0342_),
    .A4(_0409_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2132_ (.I(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2133_ (.A1(_0457_),
    .A2(_0481_),
    .B(_0483_),
    .C(_0479_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2134_ (.A1(_0343_),
    .A2(_0375_),
    .B(_0371_),
    .C(_0370_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2135_ (.A1(_0352_),
    .A2(_0375_),
    .B(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2136_ (.A1(_0484_),
    .A2(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2137_ (.A1(_0338_),
    .A2(_0388_),
    .B1(_0393_),
    .B2(_0427_),
    .C(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2138_ (.A1(_0356_),
    .A2(_0370_),
    .B1(_0393_),
    .B2(_0338_),
    .C(_0347_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2139_ (.A1(_0480_),
    .A2(_0488_),
    .B1(_0489_),
    .B2(_0345_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2140_ (.A1(_0360_),
    .A2(_0397_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _2141_ (.A1(_0360_),
    .A2(_0427_),
    .B1(_0362_),
    .B2(_0478_),
    .C1(_0491_),
    .C2(_0338_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2142_ (.A1(_0402_),
    .A2(_0492_),
    .B(_0421_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2143_ (.A1(_0405_),
    .A2(_0478_),
    .B1(_0490_),
    .B2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2144_ (.A1(_0477_),
    .A2(_0494_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2145_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_0382_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2146_ (.A1(_1016_),
    .A2(_1005_),
    .A3(_0859_),
    .B(_1029_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2147_ (.A1(_0333_),
    .A2(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2148_ (.I(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2149_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2150_ (.A1(_0495_),
    .A2(_0498_),
    .B(_0499_),
    .C(_0455_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2151_ (.I(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2152_ (.A1(_0500_),
    .A2(_0496_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2153_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_0496_),
    .B(_0501_),
    .C(_0334_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2154_ (.A1(_0464_),
    .A2(_0502_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2155_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2156_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0496_),
    .B(_0382_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2157_ (.A1(_0503_),
    .A2(_0498_),
    .B1(_0504_),
    .B2(_0476_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2158_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_0899_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2159_ (.A1(_0470_),
    .A2(_0469_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2160_ (.A1(_0343_),
    .A2(_0425_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2161_ (.A1(_0415_),
    .A2(_0507_),
    .B(_0469_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2162_ (.A1(_0427_),
    .A2(_0506_),
    .B(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2163_ (.A1(_0413_),
    .A2(_0397_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2164_ (.A1(_0385_),
    .A2(_0505_),
    .B(_0510_),
    .C(_0491_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2165_ (.A1(_0427_),
    .A2(_0433_),
    .B(_0379_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2166_ (.A1(_0379_),
    .A2(_0509_),
    .B1(_0511_),
    .B2(_0512_),
    .C(_0381_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2167_ (.A1(_0381_),
    .A2(_0505_),
    .B(_0513_),
    .C(_0382_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2168_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_1192_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2169_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0498_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2170_ (.A1(_0498_),
    .A2(_0514_),
    .A3(_0515_),
    .B(_0516_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2171_ (.A1(_0335_),
    .A2(_0388_),
    .B(_0367_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2172_ (.A1(_0350_),
    .A2(_0416_),
    .B(_0507_),
    .C(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2173_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_0900_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2174_ (.A1(_0335_),
    .A2(_0397_),
    .B1(_0401_),
    .B2(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2175_ (.A1(_0368_),
    .A2(_0350_),
    .B1(_0402_),
    .B2(_0520_),
    .C(_0403_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2176_ (.A1(_0395_),
    .A2(_0518_),
    .A3(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2177_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0333_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2178_ (.A1(_0498_),
    .A2(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2179_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_0498_),
    .B1(_0519_),
    .B2(_0405_),
    .C(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(_0522_),
    .A2(_0525_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2181_ (.A1(_0371_),
    .A2(_0375_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2182_ (.A1(_0394_),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2183_ (.A1(_0356_),
    .A2(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2184_ (.I(_0457_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2185_ (.A1(_0343_),
    .A2(_0529_),
    .B(_0482_),
    .C(_0448_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2186_ (.A1(_0345_),
    .A2(_0528_),
    .A3(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2187_ (.A1(_0343_),
    .A2(_0345_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2188_ (.A1(_0368_),
    .A2(_0399_),
    .B(_0532_),
    .C(_0381_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2189_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .S(_0900_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2190_ (.A1(_0531_),
    .A2(_0533_),
    .B1(_0534_),
    .B2(_0381_),
    .C(_0382_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2191_ (.A1(_0855_),
    .A2(_0857_),
    .A3(\u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2192_ (.A1(_1016_),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2193_ (.A1(_1029_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2194_ (.A1(_0333_),
    .A2(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2195_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_0407_),
    .B(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2196_ (.A1(_1016_),
    .A2(_0536_),
    .B(_1165_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2197_ (.A1(_1192_),
    .A2(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2198_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2199_ (.A1(_0535_),
    .A2(_0540_),
    .B(_0543_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2200_ (.A1(_1192_),
    .A2(_0538_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2201_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_0542_),
    .B1(_0544_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2202_ (.A1(_0494_),
    .A2(_0545_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2203_ (.A1(_0354_),
    .A2(_0370_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2204_ (.A1(_0426_),
    .A2(_0420_),
    .B(_0367_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2205_ (.A1(_0526_),
    .A2(_0546_),
    .B(_0547_),
    .C(_0530_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2206_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_0900_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2207_ (.A1(_0340_),
    .A2(_0433_),
    .B1(_0549_),
    .B2(_0401_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2208_ (.A1(_0340_),
    .A2(_0393_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2209_ (.A1(_0354_),
    .A2(_0370_),
    .B(_0347_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2210_ (.A1(_0402_),
    .A2(_0550_),
    .B1(_0551_),
    .B2(_0552_),
    .C(_0421_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2211_ (.A1(_0548_),
    .A2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2212_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_0542_),
    .B1(_0544_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_0549_),
    .C2(_0405_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2213_ (.A1(_0554_),
    .A2(_0555_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2214_ (.A1(_0467_),
    .A2(_0375_),
    .B(_0485_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2215_ (.A1(_0484_),
    .A2(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2216_ (.A1(_0337_),
    .A2(_0388_),
    .B1(_0393_),
    .B2(_0343_),
    .C(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2217_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .S(_0900_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2218_ (.A1(_0337_),
    .A2(_0433_),
    .B1(_0559_),
    .B2(_0401_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2219_ (.A1(_0480_),
    .A2(_0558_),
    .B1(_0560_),
    .B2(_0379_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2220_ (.A1(_0421_),
    .A2(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2221_ (.A1(_0333_),
    .A2(_0541_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2222_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_0539_),
    .B1(_0563_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2223_ (.A1(_0382_),
    .A2(_0404_),
    .A3(_0559_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2224_ (.A1(_0562_),
    .A2(_0564_),
    .A3(_0565_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2225_ (.A1(_0900_),
    .A2(\u_arbiter.i_wb_cpu_rdt[29] ),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2226_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2227_ (.A1(_0361_),
    .A2(_0567_),
    .B(_0379_),
    .C(_0385_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2228_ (.A1(_0336_),
    .A2(_0388_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2229_ (.A1(_0479_),
    .A2(_0481_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2230_ (.A1(_0482_),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2231_ (.A1(_0569_),
    .A2(_0571_),
    .B(_0480_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2232_ (.A1(_0510_),
    .A2(_0568_),
    .B(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2233_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_0539_),
    .B1(_0563_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2234_ (.A1(_0405_),
    .A2(_0567_),
    .B1(_0573_),
    .B2(_0395_),
    .C(_0574_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2235_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_0900_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2236_ (.A1(_0413_),
    .A2(_0343_),
    .B(_0411_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2237_ (.A1(_0411_),
    .A2(_0413_),
    .B1(_0442_),
    .B2(_0576_),
    .C(_0429_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2238_ (.A1(_0340_),
    .A2(_0388_),
    .B(_0570_),
    .C(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2239_ (.A1(_0480_),
    .A2(_0578_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2240_ (.A1(_0405_),
    .A2(_0575_),
    .B1(_0579_),
    .B2(_1192_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2241_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_0542_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2242_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2243_ (.A1(_0855_),
    .A2(_1016_),
    .B(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2244_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_1020_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2245_ (.A1(_0584_),
    .A2(_0583_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2246_ (.A1(_0582_),
    .A2(_0583_),
    .B(_0585_),
    .C(_1170_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2247_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_1170_),
    .B(_0544_),
    .C(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2248_ (.A1(_0580_),
    .A2(_0581_),
    .A3(_0587_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2249_ (.A1(_0339_),
    .A2(_0340_),
    .B(_0343_),
    .C(_0363_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2250_ (.A1(_0338_),
    .A2(_0398_),
    .A3(_0419_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2251_ (.A1(_0368_),
    .A2(_0588_),
    .A3(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2252_ (.A1(_0899_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2253_ (.A1(_1189_),
    .A2(\u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2254_ (.A1(_0371_),
    .A2(_0491_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2255_ (.A1(_0343_),
    .A2(_0393_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2256_ (.A1(_0592_),
    .A2(_0385_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2257_ (.A1(_0338_),
    .A2(_0409_),
    .B1(_0595_),
    .B2(_0397_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2258_ (.A1(_0592_),
    .A2(_0593_),
    .B1(_0594_),
    .B2(_0596_),
    .C(_0408_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2259_ (.A1(_0367_),
    .A2(_0590_),
    .B(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2260_ (.A1(_0397_),
    .A2(_0356_),
    .B1(_0401_),
    .B2(_0338_),
    .C(_0379_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2261_ (.A1(_0598_),
    .A2(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2262_ (.A1(_0338_),
    .A2(_0405_),
    .B1(_0600_),
    .B2(_0395_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2263_ (.A1(_1165_),
    .A2(_0584_),
    .B(_0382_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2264_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_0407_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2265_ (.A1(_0601_),
    .A2(_0602_),
    .B1(_0603_),
    .B2(_1165_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2266_ (.A1(_0856_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2267_ (.A1(_1020_),
    .A2(_1077_),
    .A3(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2268_ (.A1(_1029_),
    .A2(_0605_),
    .B(_1192_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2269_ (.I(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2270_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_0334_),
    .B(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2271_ (.A1(_0582_),
    .A2(_0607_),
    .B1(_0608_),
    .B2(_0455_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2272_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2273_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_0334_),
    .B(_0607_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2274_ (.A1(_0609_),
    .A2(_0607_),
    .B1(_0610_),
    .B2(_0436_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2275_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2276_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_0334_),
    .B(_0606_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2277_ (.A1(_0611_),
    .A2(_0607_),
    .B1(_0612_),
    .B2(_0441_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2278_ (.I(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2279_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_0334_),
    .B(_0606_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2280_ (.A1(_0613_),
    .A2(_0607_),
    .B1(_0614_),
    .B2(_0445_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2281_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2282_ (.A1(_0343_),
    .A2(_0388_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2283_ (.A1(_0352_),
    .A2(_0376_),
    .B(_0616_),
    .C(_0479_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2284_ (.A1(_0338_),
    .A2(_0479_),
    .B(_0617_),
    .C(_0369_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2285_ (.A1(_0379_),
    .A2(_0433_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2286_ (.A1(_0337_),
    .A2(_0479_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2287_ (.A1(_0408_),
    .A2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2288_ (.A1(_0397_),
    .A2(_0388_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2289_ (.A1(_0343_),
    .A2(_0397_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2290_ (.A1(_0358_),
    .A2(_0623_),
    .B(_0470_),
    .C(_0385_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2291_ (.A1(_0621_),
    .A2(_0622_),
    .B(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2292_ (.I(_0625_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2293_ (.A1(_0619_),
    .A2(_0595_),
    .B1(_0626_),
    .B2(_0338_),
    .C(_0381_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2294_ (.A1(_0397_),
    .A2(_0403_),
    .B1(_0618_),
    .B2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2295_ (.A1(_0407_),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2296_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0334_),
    .B(_0607_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2297_ (.A1(_0615_),
    .A2(_0607_),
    .B1(_0629_),
    .B2(_0630_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2298_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_0899_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2299_ (.A1(_0401_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2300_ (.A1(_0340_),
    .A2(_0385_),
    .B(_0379_),
    .C(_0433_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2301_ (.A1(_0426_),
    .A2(_0375_),
    .B(_0371_),
    .C(_0370_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(_0340_),
    .A2(_0409_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2303_ (.A1(_0616_),
    .A2(_0479_),
    .A3(_0551_),
    .A4(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2304_ (.A1(_0374_),
    .A2(_0593_),
    .B1(_0634_),
    .B2(_0636_),
    .C(_0408_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2305_ (.A1(_0358_),
    .A2(_0623_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2306_ (.A1(_0340_),
    .A2(_0348_),
    .A3(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2307_ (.A1(_0379_),
    .A2(_0399_),
    .A3(_0639_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2308_ (.A1(_0637_),
    .A2(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2309_ (.A1(_0632_),
    .A2(_0633_),
    .B(_0381_),
    .C(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2310_ (.A1(_0381_),
    .A2(_0631_),
    .B(_0642_),
    .C(_0382_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2311_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_1192_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2312_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0607_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2313_ (.A1(_0607_),
    .A2(_0643_),
    .A3(_0644_),
    .B(_0645_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2314_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .S(_0899_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2315_ (.A1(_0449_),
    .A2(_0479_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2316_ (.A1(_0337_),
    .A2(_0626_),
    .B1(_0647_),
    .B2(_0621_),
    .C(_0402_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2317_ (.A1(_0337_),
    .A2(_0385_),
    .B1(_0401_),
    .B2(_0646_),
    .C(_0379_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2318_ (.A1(_0381_),
    .A2(_0648_),
    .A3(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2319_ (.A1(_0381_),
    .A2(_0646_),
    .B(_0650_),
    .C(_0382_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2320_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_1192_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2321_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0607_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2322_ (.A1(_0607_),
    .A2(_0651_),
    .A3(_0652_),
    .B(_0653_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2323_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .S(_0900_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2324_ (.A1(_0370_),
    .A2(_0388_),
    .B(_0449_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2325_ (.A1(_0413_),
    .A2(_0593_),
    .B(_0408_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2326_ (.A1(_0336_),
    .A2(_0624_),
    .B1(_0655_),
    .B2(_0656_),
    .C(_0402_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2327_ (.A1(_0360_),
    .A2(_0402_),
    .B(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2328_ (.A1(_0381_),
    .A2(_0654_),
    .B(_0658_),
    .C(_0382_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2329_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_1192_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2330_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0607_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2331_ (.A1(_0607_),
    .A2(_0659_),
    .A3(_0660_),
    .B(_0661_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2332_ (.A1(_0411_),
    .A2(_0479_),
    .B(_0449_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2333_ (.A1(_0900_),
    .A2(_0272_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2334_ (.A1(_0900_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_0381_),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2335_ (.A1(_1192_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2336_ (.A1(_0335_),
    .A2(_0624_),
    .B1(_0662_),
    .B2(_0369_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2337_ (.A1(_0858_),
    .A2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2338_ (.A1(_0382_),
    .A2(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2339_ (.A1(_0857_),
    .A2(_0584_),
    .B(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2340_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0607_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2341_ (.A1(_0607_),
    .A2(_0666_),
    .A3(_0669_),
    .B(_0670_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2342_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_0900_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2343_ (.A1(_0616_),
    .A2(_0571_),
    .B(_0480_),
    .C(_0382_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2344_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_0334_),
    .B1(_0405_),
    .B2(_0671_),
    .C(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2345_ (.I(_0673_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2346_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2347_ (.A1(_1014_),
    .A2(_1181_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2348_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2349_ (.A1(_0674_),
    .A2(_0675_),
    .B(_0676_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2350_ (.I0(\u_cpu.cpu.alu.cmp_r ),
    .I1(_0244_),
    .S(_1029_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2351_ (.I(_0677_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2352_ (.I(_1073_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2353_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2354_ (.I(_0679_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2355_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_0678_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2356_ (.I(_0680_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2357_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_0678_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2358_ (.I(_0681_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2359_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_0678_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2360_ (.I(_0682_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2361_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_0678_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2362_ (.I(_0683_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2363_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_0678_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2364_ (.I(_0684_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2365_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_0678_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2366_ (.I(_0685_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2367_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_0678_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2368_ (.I(_0686_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2369_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_0678_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2370_ (.I(_0687_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2371_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_0678_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2372_ (.I(_0688_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2373_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_0678_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2374_ (.I(_0689_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2375_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_0678_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2376_ (.I(_0690_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2377_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_0678_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2378_ (.I(_0691_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2379_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_0678_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2380_ (.I(_0692_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2381_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_0678_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2382_ (.I(_0693_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2383_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_0678_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2384_ (.I(_0694_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2385_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_1073_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2386_ (.I(_0695_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2387_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_1073_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2388_ (.I(_0696_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2389_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_1073_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2390_ (.I(_0697_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2391_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_1073_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2392_ (.I(_0698_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2393_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_1073_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2394_ (.I(_0699_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2395_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_1073_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2396_ (.I(_0700_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2397_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_1073_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2398_ (.I(_0701_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2399_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_1073_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2400_ (.I(_0702_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2401_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_1073_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2402_ (.I(_0703_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2403_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_1073_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2404_ (.I(_0704_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2405_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_1073_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2406_ (.I(_0705_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2407_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_1073_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2408_ (.I(_0706_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2409_ (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2410_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_1064_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2411_ (.A1(_0707_),
    .A2(_1064_),
    .B(_0708_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2412_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_1181_),
    .B(_1064_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2413_ (.A1(_1173_),
    .A2(_1176_),
    .B(_1181_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2414_ (.A1(_1173_),
    .A2(_1176_),
    .B(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2415_ (.A1(_0707_),
    .A2(_0709_),
    .B1(_0711_),
    .B2(_1064_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2416_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .B(_1038_),
    .C(_1195_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2417_ (.A1(_1064_),
    .A2(_1195_),
    .B(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2418_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2419_ (.A1(_1053_),
    .A2(_0713_),
    .B(_0714_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2420_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_1181_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2421_ (.A1(_0711_),
    .A2(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2422_ (.A1(_0713_),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2423_ (.A1(_1163_),
    .A2(_0713_),
    .B(_0717_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2424_ (.A1(_1029_),
    .A2(_1181_),
    .B(_0891_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2425_ (.I(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2426_ (.A1(_0891_),
    .A2(_1182_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2427_ (.I(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2428_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2429_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2430_ (.I(_0723_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2431_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2432_ (.I(_0724_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2433_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2434_ (.I(_0725_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2435_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2436_ (.I(_0726_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2437_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2438_ (.I(_0727_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2439_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2440_ (.I(_0728_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2441_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2442_ (.I(_0729_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2443_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2444_ (.I(_0730_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2445_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2446_ (.I(_0731_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2447_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2448_ (.I(_0732_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2449_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2450_ (.I(_0733_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2451_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2452_ (.I(_0734_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2453_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2454_ (.I(_0735_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2455_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2456_ (.I(_0736_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2457_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0719_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2458_ (.I(_0737_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2459_ (.I(_0718_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2460_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_0738_),
    .B1(_0722_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2461_ (.I(_0739_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2462_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2463_ (.I(_0740_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2464_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2465_ (.I(_0741_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2466_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2467_ (.I(_0742_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2468_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2469_ (.I(_0743_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2470_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2471_ (.I(_0744_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2472_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2473_ (.I(_0745_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2474_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2475_ (.I(_0746_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2476_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2477_ (.I(_0747_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2478_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2479_ (.I(_0748_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2480_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2481_ (.I(_0749_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2482_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2483_ (.I(_0750_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2484_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2485_ (.I(_0751_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2486_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2487_ (.I(_0752_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2488_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2489_ (.I(_0753_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2490_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_0738_),
    .B1(_0721_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2491_ (.I(_0754_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2492_ (.A1(_0864_),
    .A2(_0870_),
    .A3(_0866_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2493_ (.A1(_0873_),
    .A2(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2494_ (.I(_1106_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2495_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2496_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_1081_),
    .B(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2497_ (.A1(_0756_),
    .A2(_1091_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2498_ (.A1(_0756_),
    .A2(_0759_),
    .B1(_0760_),
    .B2(_1036_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2499_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0718_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2500_ (.A1(_0891_),
    .A2(_1182_),
    .A3(_0761_),
    .B(_0762_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2501_ (.A1(_1165_),
    .A2(_1186_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2502_ (.A1(_1192_),
    .A2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2503_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0334_),
    .B(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2504_ (.A1(_1015_),
    .A2(_0764_),
    .B1(_0765_),
    .B2(_0601_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2505_ (.A1(_0340_),
    .A2(_0348_),
    .A3(_0398_),
    .A4(_0419_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2506_ (.A1(_0340_),
    .A2(_0370_),
    .B1(_0393_),
    .B2(_0354_),
    .C(_0593_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2507_ (.A1(_0374_),
    .A2(_0593_),
    .B1(_0635_),
    .B2(_0767_),
    .C(_0408_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2508_ (.A1(_0402_),
    .A2(_0768_),
    .B(_0404_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2509_ (.A1(_0397_),
    .A2(_0354_),
    .B1(_0401_),
    .B2(_0340_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2510_ (.A1(_0766_),
    .A2(_0769_),
    .B1(_0770_),
    .B2(_0402_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2511_ (.A1(_0407_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2512_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0763_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2513_ (.A1(_1159_),
    .A2(_0763_),
    .B(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2514_ (.A1(_0340_),
    .A2(_0405_),
    .B1(_0774_),
    .B2(_0334_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2515_ (.A1(_0772_),
    .A2(_0775_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2516_ (.A1(_0397_),
    .A2(_0355_),
    .B1(_0393_),
    .B2(_0426_),
    .C1(_0401_),
    .C2(_0337_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2517_ (.A1(_0337_),
    .A2(_0394_),
    .A3(_0491_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2518_ (.A1(_0473_),
    .A2(_0479_),
    .A3(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2519_ (.A1(_0621_),
    .A2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2520_ (.A1(_0379_),
    .A2(_0776_),
    .B(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2521_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0382_),
    .B1(_0395_),
    .B2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2522_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_0764_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2523_ (.A1(_0470_),
    .A2(_0363_),
    .B(_0404_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2524_ (.A1(_0407_),
    .A2(_0337_),
    .A3(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2525_ (.A1(_0764_),
    .A2(_0781_),
    .B(_0782_),
    .C(_0784_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2526_ (.A1(_1162_),
    .A2(_0763_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2527_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0763_),
    .B(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2528_ (.A1(_0368_),
    .A2(_0388_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2529_ (.A1(_0402_),
    .A2(_0783_),
    .A3(_0787_),
    .B(_0336_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2530_ (.A1(_0361_),
    .A2(_0379_),
    .B1(_0429_),
    .B2(_0408_),
    .C(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2531_ (.A1(_0407_),
    .A2(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2532_ (.A1(_0407_),
    .A2(_0786_),
    .B(_0790_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2533_ (.A1(_0345_),
    .A2(_0451_),
    .A3(_0457_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2534_ (.A1(_0398_),
    .A2(_0379_),
    .A3(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2535_ (.A1(_0404_),
    .A2(_0419_),
    .A3(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2536_ (.A1(_0382_),
    .A2(_0411_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2537_ (.A1(_0793_),
    .A2(_0794_),
    .B(_0764_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2538_ (.A1(_1162_),
    .A2(_0764_),
    .B1(_0795_),
    .B2(_0523_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2539_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_0334_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2540_ (.A1(_0580_),
    .A2(_0796_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(\u_arbiter.o_wb_cpu_adr[1] ),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2542_ (.A1(_0900_),
    .A2(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2543_ (.A1(_0891_),
    .A2(_0798_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2544_ (.I(_1190_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2545_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0799_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2546_ (.I(_0800_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2547_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_0799_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2548_ (.I(_0801_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2549_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0799_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(_0802_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2551_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_0799_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2552_ (.I(_0803_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2553_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0799_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2554_ (.I(_0804_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2555_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_0799_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2556_ (.I(_0805_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2557_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_0799_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2558_ (.I(_0806_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2559_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0799_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2560_ (.I(_0807_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2561_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_0799_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2562_ (.I(_0808_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2563_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0799_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2564_ (.I(_0809_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2565_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0799_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2566_ (.I(_0810_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2567_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0799_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2568_ (.I(_0811_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2569_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0799_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2570_ (.I(_0812_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2571_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_0799_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2572_ (.I(_0813_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2573_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0799_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2574_ (.I(_0814_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2575_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_0799_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2576_ (.I(_0815_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2577_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2578_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_0816_),
    .B(_0872_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2579_ (.A1(_1014_),
    .A2(_0873_),
    .B1(_1045_),
    .B2(_1038_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2580_ (.I0(_0817_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .S(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2581_ (.I(_0819_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2582_ (.A1(_0858_),
    .A2(\u_arbiter.i_wb_cpu_dbus_we ),
    .B1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .B2(_0869_),
    .C(_0818_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2583_ (.A1(_0816_),
    .A2(_0818_),
    .B1(_0820_),
    .B2(_0872_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2584_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2585_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2586_ (.A1(_0822_),
    .A2(_0873_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2587_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_0858_),
    .A3(_0818_),
    .A4(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2588_ (.A1(_0821_),
    .A2(_0818_),
    .B(_0824_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2589_ (.A1(_0863_),
    .A2(_0871_),
    .B(_0818_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2590_ (.A1(_0822_),
    .A2(_0818_),
    .B1(_0825_),
    .B2(_1051_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2591_ (.I(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2592_ (.A1(_1014_),
    .A2(_1044_),
    .B(_0873_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2593_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2594_ (.A1(_0826_),
    .A2(_0827_),
    .B1(_0828_),
    .B2(_1051_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2595_ (.A1(_1014_),
    .A2(_0873_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2596_ (.I0(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .I1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .S(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2597_ (.I(_0830_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2598_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2599_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .A4(_1037_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2600_ (.A1(_1039_),
    .A2(_0224_),
    .A3(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2601_ (.A1(_1050_),
    .A2(_0833_),
    .B(_0892_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2602_ (.A1(_0831_),
    .A2(_0833_),
    .B(_0834_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2603_ (.A1(_0755_),
    .A2(_1050_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2604_ (.A1(_0755_),
    .A2(_1040_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2605_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_0862_),
    .B(_0886_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2606_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_0829_),
    .A3(_0836_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2607_ (.A1(_0835_),
    .A2(_0836_),
    .A3(_0837_),
    .B(_0838_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2608_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_0334_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2609_ (.A1(_0421_),
    .A2(_0839_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2610_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_0228_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2611_ (.A1(_0891_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_0676_),
    .B(_0840_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2612_ (.A1(_0382_),
    .A2(_0228_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2613_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2614_ (.A1(_0719_),
    .A2(_0841_),
    .B(_0842_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2615_ (.A1(_1128_),
    .A2(_0024_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2616_ (.A1(_1011_),
    .A2(_0843_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2617_ (.A1(_0851_),
    .A2(_0843_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2618_ (.A1(_0892_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2619_ (.I(_0844_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2620_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0850_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(_0215_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2622_ (.A1(_0845_),
    .A2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2623_ (.A1(_1193_),
    .A2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2624_ (.A1(_1206_),
    .A2(_0848_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2625_ (.D(_0027_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2626_ (.D(_0028_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2627_ (.D(_0029_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2628_ (.D(_0030_),
    .CLK(io_in[4]),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2629_ (.D(_0031_),
    .CLK(io_in[4]),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2630_ (.D(_0007_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2631_ (.D(_0008_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2632_ (.D(_0009_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2633_ (.D(_0010_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2634_ (.D(_0011_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2635_ (.D(_0012_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2636_ (.D(_0000_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2637_ (.D(_0001_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2638_ (.D(_0002_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2639_ (.D(_0003_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2640_ (.D(_0004_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2641_ (.D(_0005_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2642_ (.D(_0006_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2643_ (.D(_0032_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2644_ (.D(_0033_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2645_ (.D(_0034_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2646_ (.D(_0035_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2647_ (.D(_0036_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2648_ (.D(_0037_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2649_ (.D(_0038_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2650_ (.D(_0039_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2651_ (.D(_0040_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2652_ (.D(_0041_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2653_ (.D(_0042_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2654_ (.D(_0043_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2655_ (.D(_0044_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2656_ (.D(_0045_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2657_ (.D(_0046_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2658_ (.D(_0047_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2659_ (.D(_0048_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2660_ (.D(_0049_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2661_ (.D(_0050_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2662_ (.D(_0051_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2663_ (.D(_0052_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2664_ (.D(_0053_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2665_ (.D(_0054_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2666_ (.D(_0055_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2667_ (.D(_0056_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2668_ (.D(_0057_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2669_ (.D(_0058_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2670_ (.D(_0059_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2671_ (.D(_0060_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2672_ (.D(_0061_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2673_ (.D(_0062_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2674_ (.D(_0063_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2675_ (.D(_0064_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2676_ (.D(_0065_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2677_ (.D(_0066_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2678_ (.D(_0067_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2679_ (.D(_0068_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2680_ (.D(_0069_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2681_ (.D(_0070_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2682_ (.D(_0071_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2683_ (.D(_0072_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2684_ (.D(_0073_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2685_ (.D(_0074_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2686_ (.D(_0075_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2687_ (.D(_0076_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2688_ (.D(_0077_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2689_ (.D(_0078_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2690_ (.D(_0079_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2691_ (.D(_0080_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2692_ (.D(_0081_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2693_ (.D(_0082_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2694_ (.D(_0083_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2695_ (.D(_0084_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2696_ (.D(_0085_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2697_ (.D(_0086_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2698_ (.D(_0087_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2699_ (.D(_0088_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2700_ (.D(_0089_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2701_ (.D(_0090_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2702_ (.D(_0091_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2703_ (.D(_0092_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2704_ (.D(_0093_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2705_ (.D(_0094_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2706_ (.D(_0095_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2707_ (.D(_0096_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2708_ (.D(_0097_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2709_ (.D(_0098_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2710_ (.D(_0099_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2711_ (.D(_0100_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2712_ (.D(_0101_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2713_ (.D(_0102_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2714_ (.D(_0103_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2715_ (.D(_0104_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2716_ (.D(_0105_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2717_ (.D(_0106_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2718_ (.D(_0107_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2719_ (.D(_0108_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2720_ (.D(_0109_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2721_ (.D(_0110_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2722_ (.D(_0111_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2723_ (.D(_0112_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2724_ (.D(_0113_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2725_ (.D(_0114_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2726_ (.D(_0115_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2727_ (.D(_0116_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2728_ (.D(_0117_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2729_ (.D(_0118_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2730_ (.D(_0119_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2731_ (.D(_0120_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2732_ (.D(_0121_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2733_ (.D(_0122_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2734_ (.D(_0123_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2735_ (.D(_0124_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2736_ (.D(_0125_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2737_ (.D(_0126_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2738_ (.D(_0127_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2739_ (.D(_0128_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2740_ (.D(_0129_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2741_ (.D(_0130_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2742_ (.D(_0131_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2743_ (.D(_0132_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2744_ (.D(_0133_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2745_ (.D(_0134_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2746_ (.D(_0135_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2747_ (.D(_0136_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2748_ (.D(_0137_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2749_ (.D(_0138_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2750_ (.D(_0139_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2751_ (.D(_0140_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2752_ (.D(_0141_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2753_ (.D(_0142_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2754_ (.D(_0014_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2755_ (.D(_0143_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2756_ (.D(_0144_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2757_ (.D(_0016_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2758_ (.D(_0015_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2759_ (.D(_0145_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2760_ (.D(_0146_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2761_ (.D(_0147_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2762_ (.D(_0148_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2763_ (.D(_0149_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2764_ (.D(_0150_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2765_ (.D(_0151_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2766_ (.D(_0152_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2767_ (.D(_0153_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2768_ (.D(_0154_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2769_ (.D(_0155_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2770_ (.D(_0156_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2771_ (.D(_0157_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2772_ (.D(_0158_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2773_ (.D(_0159_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2774_ (.D(_0160_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2775_ (.D(_0161_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2776_ (.D(_0162_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2777_ (.D(_0163_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2778_ (.D(_0164_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2779_ (.D(_0165_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2780_ (.D(_0166_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2781_ (.D(_0167_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2782_ (.D(_0168_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2783_ (.D(_0169_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2784_ (.D(_0170_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2785_ (.D(_0171_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2786_ (.D(_0172_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2787_ (.D(_0173_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2788_ (.D(_0174_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2789_ (.D(_0175_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2790_ (.D(_0176_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2791_ (.D(_0013_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2792_ (.D(_0177_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2793_ (.D(_0178_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2794_ (.D(_0179_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2795_ (.D(_0180_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2796_ (.D(_0181_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2797_ (.D(_0182_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2798_ (.D(_0183_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2799_ (.D(_0184_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2800_ (.D(_0185_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2801_ (.D(_0186_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2802_ (.D(_0187_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2803_ (.D(_0188_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2804_ (.D(_0189_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2805_ (.D(_0190_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2806_ (.D(_0191_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2807_ (.D(_0192_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2808_ (.D(_0193_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2809_ (.D(_0194_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2810_ (.D(_0195_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2811_ (.D(_0196_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2812_ (.D(_0197_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2813_ (.D(_0198_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2814_ (.D(_0199_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2815_ (.D(_0200_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2816_ (.D(_0201_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2817_ (.D(_0202_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2818_ (.D(_0203_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2819_ (.D(_0204_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2820_ (.D(_0205_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2821_ (.D(_0206_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2822_ (.D(_0207_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2823_ (.D(_0208_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2824_ (.D(_0209_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2825_ (.D(_0017_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2826_ (.D(_0018_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2827_ (.D(_0019_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2828_ (.D(_0020_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2829_ (.D(_0021_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2830_ (.D(_0022_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2831_ (.D(_0023_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2832_ (.D(_0024_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2833_ (.D(_0025_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2834_ (.D(_0210_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2835_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2836_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2837_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2838_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2839_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2840_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2841_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2842_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2843_ (.D(_0211_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2844_ (.D(_0212_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2845_ (.D(_0213_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2846_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2847_ (.D(_0214_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2848_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2849_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2850_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2851_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2852_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2853_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2854_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2855_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2856_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2857_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2858_ (.Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2859_ (.Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2860_ (.Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2861_ (.Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2862_ (.Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2863_ (.Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2864_ (.Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2865_ (.Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2866_ (.Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2867_ (.Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2868_ (.Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2869_ (.Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2870_ (.Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2871_ (.Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2872_ (.Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2873_ (.Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2874_ (.Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2875_ (.Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2876_ (.Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2877_ (.Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2878_ (.Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2879_ (.Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2880_ (.Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2881_ (.Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2882_ (.Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2883_ (.Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2884_ (.Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2885_ (.Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2886_ (.Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2887_ (.Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2888_ (.Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2889_ (.Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2890_ (.Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2891_ (.Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2892_ (.Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2893_ (.Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2894_ (.Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2895_ (.Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2896_ (.Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2897_ (.Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2898_ (.Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2899_ (.Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2900_ (.Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2901_ (.Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2902_ (.Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2903_ (.Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2904_ (.Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2905_ (.Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2906_ (.Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2907_ (.Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2908_ (.Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2909_ (.Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2910_ (.Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2911_ (.Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2912_ (.Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2913_ (.Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2914_ (.Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2915_ (.Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2916_ (.Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2917_ (.Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2918_ (.Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2919_ (.Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2920_ (.Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2921_ (.Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2922_ (.Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2923_ (.Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2924_ (.Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2925_ (.Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2926_ (.Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2927_ (.Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2928_ (.Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2929_ (.Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2930_ (.Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2931_ (.Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2932_ (.ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2933_ (.ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2934_ (.ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2935_ (.ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2936_ (.ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2937_ (.ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2938_ (.ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2939_ (.ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2940_ (.ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2941_ (.ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2942_ (.ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2943_ (.ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2944_ (.ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2945_ (.ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2946_ (.ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2947_ (.ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2948_ (.ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2949_ (.ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2950_ (.ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2951_ (.ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2952_ (.ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2953_ (.ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2954_ (.ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2955_ (.ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2956_ (.ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2957_ (.ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2958_ (.ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2959_ (.ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2960_ (.ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2961_ (.ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2962_ (.ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2963_ (.ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2964_ (.ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2965_ (.ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2966_ (.ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2967_ (.ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2968_ (.ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2969_ (.ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2970_ (.ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2971_ (.ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2972_ (.ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2973_ (.ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2974_ (.ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2975_ (.ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2976_ (.ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2977_ (.ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2978_ (.ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2979_ (.ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2980_ (.ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2981_ (.ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2982_ (.ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2983_ (.ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2984_ (.ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2985_ (.ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2986_ (.ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2987_ (.ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2988_ (.ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2989_ (.ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2990_ (.ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2991_ (.ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2992_ (.ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2993_ (.ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2994_ (.ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2995_ (.ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2996_ (.ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2997_ (.ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2998_ (.ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2999_ (.ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3000_ (.ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3001_ (.ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3002_ (.ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3003_ (.ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3004_ (.ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3005_ (.ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3006_ (.ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3007_ (.ZN(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3008_ (.ZN(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3009_ (.ZN(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3010_ (.ZN(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3011_ (.ZN(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3012_ (.ZN(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3013_ (.ZN(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3014_ (.ZN(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3015_ (.I(\u_scanchain_local.clk_out ),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3016_ (.I(\u_scanchain_local.data_out ),
    .Z(io_out[1]));
 gf180mcu_fd_ip_sram__sram256x8m8wm1 \u_cpu.rf_ram.RAM0  (.CEN(_1282_),
    .CLK(io_in[4]),
    .GWEN(_0026_),
    .A({\u_cpu.rf_ram.addr[7] ,
    \u_cpu.rf_ram.addr[6] ,
    \u_cpu.rf_ram.addr[5] ,
    \u_cpu.rf_ram.addr[4] ,
    \u_cpu.rf_ram.addr[3] ,
    \u_cpu.rf_ram.addr[2] ,
    \u_cpu.rf_ram.addr[1] ,
    \u_cpu.rf_ram.addr[0] }),
    .D({\u_cpu.rf_ram.i_wdata[7] ,
    \u_cpu.rf_ram.i_wdata[6] ,
    \u_cpu.rf_ram.i_wdata[5] ,
    \u_cpu.rf_ram.i_wdata[4] ,
    \u_cpu.rf_ram.i_wdata[3] ,
    \u_cpu.rf_ram.i_wdata[2] ,
    \u_cpu.rf_ram.i_wdata[1] ,
    \u_cpu.rf_ram.i_wdata[0] }),
    .Q({\u_cpu.rf_ram.data[7] ,
    \u_cpu.rf_ram.data[6] ,
    \u_cpu.rf_ram.data[5] ,
    \u_cpu.rf_ram.data[4] ,
    \u_cpu.rf_ram.data[3] ,
    \u_cpu.rf_ram.data[2] ,
    \u_cpu.rf_ram.data[1] ,
    \u_cpu.rf_ram.data[0] }),
    .WEN({_0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_}));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \u_scanchain_local.input_buf_clk  (.I(io_in[0]),
    .Z(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 \u_scanchain_local.out_flop  (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \u_scanchain_local.output_buffers[2]  (.I(\u_scanchain_local.data_out_i ),
    .Z(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \u_scanchain_local.output_buffers[3]  (.I(\u_scanchain_local.clk ),
    .Z(\u_scanchain_local.clk_out ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[0]  (.D(io_in[2]),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_cyc ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[10]  (.D(\u_arbiter.i_wb_cpu_rdt[7] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[11]  (.D(\u_arbiter.i_wb_cpu_rdt[8] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[12]  (.D(\u_arbiter.i_wb_cpu_rdt[9] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[13]  (.D(\u_arbiter.i_wb_cpu_rdt[10] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[14]  (.D(\u_arbiter.i_wb_cpu_rdt[11] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[15]  (.D(\u_arbiter.i_wb_cpu_rdt[12] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[16]  (.D(\u_arbiter.i_wb_cpu_rdt[13] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[17]  (.D(\u_arbiter.i_wb_cpu_rdt[14] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[18]  (.D(\u_arbiter.i_wb_cpu_rdt[15] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[19]  (.D(\u_arbiter.i_wb_cpu_rdt[16] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[1]  (.D(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_we ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[20]  (.D(\u_arbiter.i_wb_cpu_rdt[17] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[21]  (.D(\u_arbiter.i_wb_cpu_rdt[18] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[22]  (.D(\u_arbiter.i_wb_cpu_rdt[19] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[23]  (.D(\u_arbiter.i_wb_cpu_rdt[20] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[24]  (.D(\u_arbiter.i_wb_cpu_rdt[21] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[25]  (.D(\u_arbiter.i_wb_cpu_rdt[22] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[26]  (.D(\u_arbiter.i_wb_cpu_rdt[23] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[27]  (.D(\u_arbiter.i_wb_cpu_rdt[24] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[28]  (.D(\u_arbiter.i_wb_cpu_rdt[25] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[29]  (.D(\u_arbiter.i_wb_cpu_rdt[26] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[2]  (.D(\u_arbiter.i_wb_cpu_ack ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[0] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[30]  (.D(\u_arbiter.i_wb_cpu_rdt[27] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[31]  (.D(\u_arbiter.i_wb_cpu_rdt[28] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[32]  (.D(\u_arbiter.i_wb_cpu_rdt[29] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[33]  (.D(\u_arbiter.i_wb_cpu_rdt[30] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[34]  (.D(\u_arbiter.i_wb_cpu_rdt[31] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[35]  (.D(\u_scanchain_local.module_data_in[34] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[36]  (.D(\u_scanchain_local.module_data_in[35] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[37]  (.D(\u_scanchain_local.module_data_in[36] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[38]  (.D(\u_scanchain_local.module_data_in[37] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[0] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[39]  (.D(\u_scanchain_local.module_data_in[38] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[1] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[3]  (.D(\u_arbiter.i_wb_cpu_rdt[0] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[1] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[40]  (.D(\u_scanchain_local.module_data_in[39] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[2] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[41]  (.D(\u_scanchain_local.module_data_in[40] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[3] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[42]  (.D(\u_scanchain_local.module_data_in[41] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[4] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[43]  (.D(\u_scanchain_local.module_data_in[42] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[5] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[44]  (.D(\u_scanchain_local.module_data_in[43] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[6] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[45]  (.D(\u_scanchain_local.module_data_in[44] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[7] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[46]  (.D(\u_scanchain_local.module_data_in[45] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[8] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[47]  (.D(\u_scanchain_local.module_data_in[46] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[9] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[48]  (.D(\u_scanchain_local.module_data_in[47] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[10] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[49]  (.D(\u_scanchain_local.module_data_in[48] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[11] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[4]  (.D(\u_arbiter.i_wb_cpu_rdt[1] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[2] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[50]  (.D(\u_scanchain_local.module_data_in[49] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[12] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[51]  (.D(\u_scanchain_local.module_data_in[50] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[13] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[52]  (.D(\u_scanchain_local.module_data_in[51] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[14] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[53]  (.D(\u_scanchain_local.module_data_in[52] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[15] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[54]  (.D(\u_scanchain_local.module_data_in[53] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[16] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[55]  (.D(\u_scanchain_local.module_data_in[54] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[17] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[56]  (.D(\u_scanchain_local.module_data_in[55] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[18] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[57]  (.D(\u_scanchain_local.module_data_in[56] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[19] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[58]  (.D(\u_scanchain_local.module_data_in[57] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[20] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[59]  (.D(\u_scanchain_local.module_data_in[58] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[21] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[5]  (.D(\u_arbiter.i_wb_cpu_rdt[2] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[3] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[60]  (.D(\u_scanchain_local.module_data_in[59] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[22] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[61]  (.D(\u_scanchain_local.module_data_in[60] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[23] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[62]  (.D(\u_scanchain_local.module_data_in[61] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[24] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[63]  (.D(\u_scanchain_local.module_data_in[62] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[25] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[64]  (.D(\u_scanchain_local.module_data_in[63] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[26] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[65]  (.D(\u_scanchain_local.module_data_in[64] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[27] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[66]  (.D(\u_scanchain_local.module_data_in[65] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[28] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[67]  (.D(\u_scanchain_local.module_data_in[66] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[29] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[68]  (.D(\u_scanchain_local.module_data_in[67] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[30] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[69]  (.D(\u_scanchain_local.module_data_in[68] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[31] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[6]  (.D(\u_arbiter.i_wb_cpu_rdt[3] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[7]  (.D(\u_arbiter.i_wb_cpu_rdt[4] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[8]  (.D(\u_arbiter.i_wb_cpu_rdt[5] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[9]  (.D(\u_arbiter.i_wb_cpu_rdt[6] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__D (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A2 (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__D (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__D (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A2 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__B (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A2 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A2 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[0]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[1]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[2]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[3]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[5]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[4]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_GWEN  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[6]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[7]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A3 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__B (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__B (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__I (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__B1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__B1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A2 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__C1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__I (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__B1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__C (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__B1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__B1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__B1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__B1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__C (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__B (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__C2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A3 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__B2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__B2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__C2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__B2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A4 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__B (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__B2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__B2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__B (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__C (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__C (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__B2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__B2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__B2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__B2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__B2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A3 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__C (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__C (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__B2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__C (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__B (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__B (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__C (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__C (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__B2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__C (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__B (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__C (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__B (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__B2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__B (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__C (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__B (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__B (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__B (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__C (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__B2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__C (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__C (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__B2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__B1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__B (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__B (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__C (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__C (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__C (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__B1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__B1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__B1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__B1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__B1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__B1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__B1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__B2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__B2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__B2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__B (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__B2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__B (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__B (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__C1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__B1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__B1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__B2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__B1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__B1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__C (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__C (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__B1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__C (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__C2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__B2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__B1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__B2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__B2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__C (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__B (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__C (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__C (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__B2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A4 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__B1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__B1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__B (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__B (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__B (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A4 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A3 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A3 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__C (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__B2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__B2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__B1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__C (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__B (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__C (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__B1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__B2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__B2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__B (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__C (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__B (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__B (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__B (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A3 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__B2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__C (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__B (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A3 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__B (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__B2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__B2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__B (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__B2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__C (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__C (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__B (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__I (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A3 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__C (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__C1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__B (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__B1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__B2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__B1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__C1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__B1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A3 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A3 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__C (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__B1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__B (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__B2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__B (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__B2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__B (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A3 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A3 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A3 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__S (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__B (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A3 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__C (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__S (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__B (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1395__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1387__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__C (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__S0 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__I (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A3 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1364__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__B (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__B (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__C (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__C (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__C (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A3 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__C (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__B (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__B1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__B2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__A4 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1385__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__B1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1378__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A3 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A4 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1381__A3 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__B (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A3 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__C (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__B2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__B (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__B (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__S (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__S (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1436__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1417__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__S (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__S (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__S (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__S (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__I (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__S (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__S (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__S (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__S (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__S (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__S (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1414__I (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__S (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__B (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__B (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1424__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__B (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1433__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1429__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__A4 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1435__A3 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1496__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A3 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A3 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1466__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A3 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A4 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A3 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A3 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__A4 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A3 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A3 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__S (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A3 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__B (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__I (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__S (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__S (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__S (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__S (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__S (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__S (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__I (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A3 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__I (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__C (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__B (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__B2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A3 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A3 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__S (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__B (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__S (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__B (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__B (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__B (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__B2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A4 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__B2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__B (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A3 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A4 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__B (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__B1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__B2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__B (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__B (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__S (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__I (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__I0 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__B (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A4 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__I (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__I (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__B2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__B2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__B2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A3 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__B (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__C (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__B (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__B (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__B2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__C (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__B (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__C (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__B (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__B (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__B (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__B2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A3 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A4 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_CEN  (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.input_buf_clk_I  (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_D  (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[50]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[51]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[52]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[58]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_CLK  (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_D  (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__I (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__I0 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A4 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A2 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A3 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A2 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A2 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__I (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__B (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__B2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_D  (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_D  (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A2 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_D  (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_D  (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_D  (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_D  (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_D  (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_D  (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_D  (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_D  (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_D  (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A1 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_D  (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__I0 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A2 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_D  (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_D  (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_D  (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_D  (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_D  (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_D  (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_D  (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_D  (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_D  (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_D  (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_D  (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__I1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__I0 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_D  (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_D  (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_D  (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A2 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_D  (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_D  (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A2 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_D  (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_D  (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_D  (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__I1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__I (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__I (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__B (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__I (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__S1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__A2 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__I (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A2 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A3 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__A3 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1539__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__I (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A2 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__B (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__A1 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A3 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__I0 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__B2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A4 (.I(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A1 (.I(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__I (.I(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A3 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1387__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__B2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__B2 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__B (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__B1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__D (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__I1 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A2 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__A2 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__I (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__C (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A2 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A1 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A1 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__I (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A1 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A3 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A3 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[0]  (.I(\u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[1]  (.I(\u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[2]  (.I(\u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[3]  (.I(\u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[4]  (.I(\u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[5]  (.I(\u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[6]  (.I(\u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[7]  (.I(\u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(\u_cpu.rf_ram.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__I1 (.I(\u_cpu.rf_ram.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__I1 (.I(\u_cpu.rf_ram.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__I1 (.I(\u_cpu.rf_ram.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__I1 (.I(\u_cpu.rf_ram.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__I1 (.I(\u_cpu.rf_ram.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__I1 (.I(\u_cpu.rf_ram.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__I1 (.I(\u_cpu.rf_ram.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[0]  (.I(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[1]  (.I(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[2]  (.I(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[3]  (.I(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[4]  (.I(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[5]  (.I(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[6]  (.I(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[7]  (.I(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1388__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__D (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__D (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__D (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__D (.I(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__D (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__I0 (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[51]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[52]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[50]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_CLKN  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[58]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.output_buffers[3]_I  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_D  (.I(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
endmodule

