magic
tech gf180mcuC
magscale 1 5
timestamp 1670028288
<< obsm1 >>
rect 672 855 68320 78497
<< metal2 >>
rect 336 79600 392 79900
rect 1008 79600 1064 79900
rect 1680 79600 1736 79900
rect 2352 79600 2408 79900
rect 3024 79600 3080 79900
rect 3696 79600 3752 79900
rect 4368 79600 4424 79900
rect 5376 79600 5432 79900
rect 6048 79600 6104 79900
rect 6720 79600 6776 79900
rect 7392 79600 7448 79900
rect 8064 79600 8120 79900
rect 8736 79600 8792 79900
rect 9408 79600 9464 79900
rect 10080 79600 10136 79900
rect 11088 79600 11144 79900
rect 11760 79600 11816 79900
rect 12432 79600 12488 79900
rect 13104 79600 13160 79900
rect 13776 79600 13832 79900
rect 14448 79600 14504 79900
rect 15120 79600 15176 79900
rect 16128 79600 16184 79900
rect 16800 79600 16856 79900
rect 17472 79600 17528 79900
rect 18144 79600 18200 79900
rect 18816 79600 18872 79900
rect 19488 79600 19544 79900
rect 20160 79600 20216 79900
rect 20832 79600 20888 79900
rect 21840 79600 21896 79900
rect 22512 79600 22568 79900
rect 23184 79600 23240 79900
rect 23856 79600 23912 79900
rect 24528 79600 24584 79900
rect 25200 79600 25256 79900
rect 25872 79600 25928 79900
rect 26880 79600 26936 79900
rect 27552 79600 27608 79900
rect 28224 79600 28280 79900
rect 28896 79600 28952 79900
rect 29568 79600 29624 79900
rect 30240 79600 30296 79900
rect 30912 79600 30968 79900
rect 31584 79600 31640 79900
rect 32592 79600 32648 79900
rect 33264 79600 33320 79900
rect 33936 79600 33992 79900
rect 34608 79600 34664 79900
rect 35280 79600 35336 79900
rect 35952 79600 36008 79900
rect 36624 79600 36680 79900
rect 37632 79600 37688 79900
rect 38304 79600 38360 79900
rect 38976 79600 39032 79900
rect 39648 79600 39704 79900
rect 40320 79600 40376 79900
rect 40992 79600 41048 79900
rect 41664 79600 41720 79900
rect 42672 79600 42728 79900
rect 43344 79600 43400 79900
rect 44016 79600 44072 79900
rect 44688 79600 44744 79900
rect 45360 79600 45416 79900
rect 46032 79600 46088 79900
rect 46704 79600 46760 79900
rect 47376 79600 47432 79900
rect 48384 79600 48440 79900
rect 49056 79600 49112 79900
rect 49728 79600 49784 79900
rect 50400 79600 50456 79900
rect 51072 79600 51128 79900
rect 51744 79600 51800 79900
rect 52416 79600 52472 79900
rect 53424 79600 53480 79900
rect 54096 79600 54152 79900
rect 54768 79600 54824 79900
rect 55440 79600 55496 79900
rect 56112 79600 56168 79900
rect 56784 79600 56840 79900
rect 57456 79600 57512 79900
rect 58128 79600 58184 79900
rect 59136 79600 59192 79900
rect 59808 79600 59864 79900
rect 60480 79600 60536 79900
rect 61152 79600 61208 79900
rect 61824 79600 61880 79900
rect 62496 79600 62552 79900
rect 63168 79600 63224 79900
rect 64176 79600 64232 79900
rect 64848 79600 64904 79900
rect 65520 79600 65576 79900
rect 66192 79600 66248 79900
rect 66864 79600 66920 79900
rect 67536 79600 67592 79900
rect 68208 79600 68264 79900
rect 68880 79600 68936 79900
rect 0 100 56 400
rect 672 100 728 400
rect 1344 100 1400 400
rect 2016 100 2072 400
rect 2688 100 2744 400
rect 3360 100 3416 400
rect 4032 100 4088 400
rect 4704 100 4760 400
rect 5712 100 5768 400
rect 6384 100 6440 400
rect 7056 100 7112 400
rect 7728 100 7784 400
rect 8400 100 8456 400
rect 9072 100 9128 400
rect 9744 100 9800 400
rect 10752 100 10808 400
rect 11424 100 11480 400
rect 12096 100 12152 400
rect 12768 100 12824 400
rect 13440 100 13496 400
rect 14112 100 14168 400
rect 14784 100 14840 400
rect 15456 100 15512 400
rect 16464 100 16520 400
rect 17136 100 17192 400
rect 17808 100 17864 400
rect 18480 100 18536 400
rect 19152 100 19208 400
rect 19824 100 19880 400
rect 20496 100 20552 400
rect 21504 100 21560 400
rect 22176 100 22232 400
rect 22848 100 22904 400
rect 23520 100 23576 400
rect 24192 100 24248 400
rect 24864 100 24920 400
rect 25536 100 25592 400
rect 26208 100 26264 400
rect 27216 100 27272 400
rect 27888 100 27944 400
rect 28560 100 28616 400
rect 29232 100 29288 400
rect 29904 100 29960 400
rect 30576 100 30632 400
rect 31248 100 31304 400
rect 32256 100 32312 400
rect 32928 100 32984 400
rect 33600 100 33656 400
rect 34272 100 34328 400
rect 34944 100 35000 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 37296 100 37352 400
rect 37968 100 38024 400
rect 38640 100 38696 400
rect 39312 100 39368 400
rect 39984 100 40040 400
rect 40656 100 40712 400
rect 41328 100 41384 400
rect 42000 100 42056 400
rect 43008 100 43064 400
rect 43680 100 43736 400
rect 44352 100 44408 400
rect 45024 100 45080 400
rect 45696 100 45752 400
rect 46368 100 46424 400
rect 47040 100 47096 400
rect 48048 100 48104 400
rect 48720 100 48776 400
rect 49392 100 49448 400
rect 50064 100 50120 400
rect 50736 100 50792 400
rect 51408 100 51464 400
rect 52080 100 52136 400
rect 52752 100 52808 400
rect 53760 100 53816 400
rect 54432 100 54488 400
rect 55104 100 55160 400
rect 55776 100 55832 400
rect 56448 100 56504 400
rect 57120 100 57176 400
rect 57792 100 57848 400
rect 58800 100 58856 400
rect 59472 100 59528 400
rect 60144 100 60200 400
rect 60816 100 60872 400
rect 61488 100 61544 400
rect 62160 100 62216 400
rect 62832 100 62888 400
rect 63504 100 63560 400
rect 64512 100 64568 400
rect 65184 100 65240 400
rect 65856 100 65912 400
rect 66528 100 66584 400
rect 67200 100 67256 400
rect 67872 100 67928 400
rect 68544 100 68600 400
<< obsm2 >>
rect 14 79570 306 79600
rect 422 79570 978 79600
rect 1094 79570 1650 79600
rect 1766 79570 2322 79600
rect 2438 79570 2994 79600
rect 3110 79570 3666 79600
rect 3782 79570 4338 79600
rect 4454 79570 5346 79600
rect 5462 79570 6018 79600
rect 6134 79570 6690 79600
rect 6806 79570 7362 79600
rect 7478 79570 8034 79600
rect 8150 79570 8706 79600
rect 8822 79570 9378 79600
rect 9494 79570 10050 79600
rect 10166 79570 11058 79600
rect 11174 79570 11730 79600
rect 11846 79570 12402 79600
rect 12518 79570 13074 79600
rect 13190 79570 13746 79600
rect 13862 79570 14418 79600
rect 14534 79570 15090 79600
rect 15206 79570 16098 79600
rect 16214 79570 16770 79600
rect 16886 79570 17442 79600
rect 17558 79570 18114 79600
rect 18230 79570 18786 79600
rect 18902 79570 19458 79600
rect 19574 79570 20130 79600
rect 20246 79570 20802 79600
rect 20918 79570 21810 79600
rect 21926 79570 22482 79600
rect 22598 79570 23154 79600
rect 23270 79570 23826 79600
rect 23942 79570 24498 79600
rect 24614 79570 25170 79600
rect 25286 79570 25842 79600
rect 25958 79570 26850 79600
rect 26966 79570 27522 79600
rect 27638 79570 28194 79600
rect 28310 79570 28866 79600
rect 28982 79570 29538 79600
rect 29654 79570 30210 79600
rect 30326 79570 30882 79600
rect 30998 79570 31554 79600
rect 31670 79570 32562 79600
rect 32678 79570 33234 79600
rect 33350 79570 33906 79600
rect 34022 79570 34578 79600
rect 34694 79570 35250 79600
rect 35366 79570 35922 79600
rect 36038 79570 36594 79600
rect 36710 79570 37602 79600
rect 37718 79570 38274 79600
rect 38390 79570 38946 79600
rect 39062 79570 39618 79600
rect 39734 79570 40290 79600
rect 40406 79570 40962 79600
rect 41078 79570 41634 79600
rect 41750 79570 42642 79600
rect 42758 79570 43314 79600
rect 43430 79570 43986 79600
rect 44102 79570 44658 79600
rect 44774 79570 45330 79600
rect 45446 79570 46002 79600
rect 46118 79570 46674 79600
rect 46790 79570 47346 79600
rect 47462 79570 48354 79600
rect 48470 79570 49026 79600
rect 49142 79570 49698 79600
rect 49814 79570 50370 79600
rect 50486 79570 51042 79600
rect 51158 79570 51714 79600
rect 51830 79570 52386 79600
rect 52502 79570 53394 79600
rect 53510 79570 54066 79600
rect 54182 79570 54738 79600
rect 54854 79570 55410 79600
rect 55526 79570 56082 79600
rect 56198 79570 56754 79600
rect 56870 79570 57426 79600
rect 57542 79570 58098 79600
rect 58214 79570 59106 79600
rect 59222 79570 59778 79600
rect 59894 79570 60450 79600
rect 60566 79570 61122 79600
rect 61238 79570 61794 79600
rect 61910 79570 62466 79600
rect 62582 79570 63138 79600
rect 63254 79570 64146 79600
rect 64262 79570 64818 79600
rect 64934 79570 65490 79600
rect 65606 79570 66162 79600
rect 66278 79570 66834 79600
rect 66950 79570 67506 79600
rect 67622 79570 68178 79600
rect 68294 79570 68642 79600
rect 14 430 68642 79570
rect 86 400 642 430
rect 758 400 1314 430
rect 1430 400 1986 430
rect 2102 400 2658 430
rect 2774 400 3330 430
rect 3446 400 4002 430
rect 4118 400 4674 430
rect 4790 400 5682 430
rect 5798 400 6354 430
rect 6470 400 7026 430
rect 7142 400 7698 430
rect 7814 400 8370 430
rect 8486 400 9042 430
rect 9158 400 9714 430
rect 9830 400 10722 430
rect 10838 400 11394 430
rect 11510 400 12066 430
rect 12182 400 12738 430
rect 12854 400 13410 430
rect 13526 400 14082 430
rect 14198 400 14754 430
rect 14870 400 15426 430
rect 15542 400 16434 430
rect 16550 400 17106 430
rect 17222 400 17778 430
rect 17894 400 18450 430
rect 18566 400 19122 430
rect 19238 400 19794 430
rect 19910 400 20466 430
rect 20582 400 21474 430
rect 21590 400 22146 430
rect 22262 400 22818 430
rect 22934 400 23490 430
rect 23606 400 24162 430
rect 24278 400 24834 430
rect 24950 400 25506 430
rect 25622 400 26178 430
rect 26294 400 27186 430
rect 27302 400 27858 430
rect 27974 400 28530 430
rect 28646 400 29202 430
rect 29318 400 29874 430
rect 29990 400 30546 430
rect 30662 400 31218 430
rect 31334 400 32226 430
rect 32342 400 32898 430
rect 33014 400 33570 430
rect 33686 400 34242 430
rect 34358 400 34914 430
rect 35030 400 35586 430
rect 35702 400 36258 430
rect 36374 400 37266 430
rect 37382 400 37938 430
rect 38054 400 38610 430
rect 38726 400 39282 430
rect 39398 400 39954 430
rect 40070 400 40626 430
rect 40742 400 41298 430
rect 41414 400 41970 430
rect 42086 400 42978 430
rect 43094 400 43650 430
rect 43766 400 44322 430
rect 44438 400 44994 430
rect 45110 400 45666 430
rect 45782 400 46338 430
rect 46454 400 47010 430
rect 47126 400 48018 430
rect 48134 400 48690 430
rect 48806 400 49362 430
rect 49478 400 50034 430
rect 50150 400 50706 430
rect 50822 400 51378 430
rect 51494 400 52050 430
rect 52166 400 52722 430
rect 52838 400 53730 430
rect 53846 400 54402 430
rect 54518 400 55074 430
rect 55190 400 55746 430
rect 55862 400 56418 430
rect 56534 400 57090 430
rect 57206 400 57762 430
rect 57878 400 58770 430
rect 58886 400 59442 430
rect 59558 400 60114 430
rect 60230 400 60786 430
rect 60902 400 61458 430
rect 61574 400 62130 430
rect 62246 400 62802 430
rect 62918 400 63474 430
rect 63590 400 64482 430
rect 64598 400 65154 430
rect 65270 400 65826 430
rect 65942 400 66498 430
rect 66614 400 67170 430
rect 67286 400 67842 430
rect 67958 400 68514 430
rect 68630 400 68642 430
<< metal3 >>
rect 100 79296 400 79352
rect 68600 78960 68900 79016
rect 100 78624 400 78680
rect 68600 78288 68900 78344
rect 100 77952 400 78008
rect 68600 77616 68900 77672
rect 100 77280 400 77336
rect 68600 76944 68900 77000
rect 100 76608 400 76664
rect 68600 76272 68900 76328
rect 100 75936 400 75992
rect 68600 75600 68900 75656
rect 100 75264 400 75320
rect 68600 74928 68900 74984
rect 100 74256 400 74312
rect 68600 73920 68900 73976
rect 100 73584 400 73640
rect 68600 73248 68900 73304
rect 100 72912 400 72968
rect 68600 72576 68900 72632
rect 100 72240 400 72296
rect 68600 71904 68900 71960
rect 100 71568 400 71624
rect 68600 71232 68900 71288
rect 100 70896 400 70952
rect 68600 70560 68900 70616
rect 100 70224 400 70280
rect 68600 69888 68900 69944
rect 100 69552 400 69608
rect 68600 68880 68900 68936
rect 100 68544 400 68600
rect 68600 68208 68900 68264
rect 100 67872 400 67928
rect 68600 67536 68900 67592
rect 100 67200 400 67256
rect 68600 66864 68900 66920
rect 100 66528 400 66584
rect 68600 66192 68900 66248
rect 100 65856 400 65912
rect 68600 65520 68900 65576
rect 100 65184 400 65240
rect 68600 64848 68900 64904
rect 100 64512 400 64568
rect 68600 64176 68900 64232
rect 100 63504 400 63560
rect 68600 63168 68900 63224
rect 100 62832 400 62888
rect 68600 62496 68900 62552
rect 100 62160 400 62216
rect 68600 61824 68900 61880
rect 100 61488 400 61544
rect 68600 61152 68900 61208
rect 100 60816 400 60872
rect 68600 60480 68900 60536
rect 100 60144 400 60200
rect 68600 59808 68900 59864
rect 100 59472 400 59528
rect 68600 59136 68900 59192
rect 100 58800 400 58856
rect 68600 58128 68900 58184
rect 100 57792 400 57848
rect 68600 57456 68900 57512
rect 100 57120 400 57176
rect 68600 56784 68900 56840
rect 100 56448 400 56504
rect 68600 56112 68900 56168
rect 100 55776 400 55832
rect 68600 55440 68900 55496
rect 100 55104 400 55160
rect 68600 54768 68900 54824
rect 100 54432 400 54488
rect 68600 54096 68900 54152
rect 100 53760 400 53816
rect 68600 53424 68900 53480
rect 100 52752 400 52808
rect 68600 52416 68900 52472
rect 100 52080 400 52136
rect 68600 51744 68900 51800
rect 100 51408 400 51464
rect 68600 51072 68900 51128
rect 100 50736 400 50792
rect 68600 50400 68900 50456
rect 100 50064 400 50120
rect 68600 49728 68900 49784
rect 100 49392 400 49448
rect 68600 49056 68900 49112
rect 100 48720 400 48776
rect 68600 48384 68900 48440
rect 100 48048 400 48104
rect 68600 47376 68900 47432
rect 100 47040 400 47096
rect 68600 46704 68900 46760
rect 100 46368 400 46424
rect 68600 46032 68900 46088
rect 100 45696 400 45752
rect 68600 45360 68900 45416
rect 100 45024 400 45080
rect 68600 44688 68900 44744
rect 100 44352 400 44408
rect 68600 44016 68900 44072
rect 100 43680 400 43736
rect 68600 43344 68900 43400
rect 100 43008 400 43064
rect 68600 42672 68900 42728
rect 100 42000 400 42056
rect 68600 41664 68900 41720
rect 100 41328 400 41384
rect 68600 40992 68900 41048
rect 100 40656 400 40712
rect 68600 40320 68900 40376
rect 100 39984 400 40040
rect 68600 39648 68900 39704
rect 100 39312 400 39368
rect 68600 38976 68900 39032
rect 100 38640 400 38696
rect 68600 38304 68900 38360
rect 100 37968 400 38024
rect 68600 37632 68900 37688
rect 100 36960 400 37016
rect 68600 36624 68900 36680
rect 100 36288 400 36344
rect 68600 35952 68900 36008
rect 100 35616 400 35672
rect 68600 35280 68900 35336
rect 100 34944 400 35000
rect 68600 34608 68900 34664
rect 100 34272 400 34328
rect 68600 33936 68900 33992
rect 100 33600 400 33656
rect 68600 33264 68900 33320
rect 100 32928 400 32984
rect 68600 32592 68900 32648
rect 100 32256 400 32312
rect 68600 31584 68900 31640
rect 100 31248 400 31304
rect 68600 30912 68900 30968
rect 100 30576 400 30632
rect 68600 30240 68900 30296
rect 100 29904 400 29960
rect 68600 29568 68900 29624
rect 100 29232 400 29288
rect 68600 28896 68900 28952
rect 100 28560 400 28616
rect 68600 28224 68900 28280
rect 100 27888 400 27944
rect 68600 27552 68900 27608
rect 100 27216 400 27272
rect 68600 26880 68900 26936
rect 100 26208 400 26264
rect 68600 25872 68900 25928
rect 100 25536 400 25592
rect 68600 25200 68900 25256
rect 100 24864 400 24920
rect 68600 24528 68900 24584
rect 100 24192 400 24248
rect 68600 23856 68900 23912
rect 100 23520 400 23576
rect 68600 23184 68900 23240
rect 100 22848 400 22904
rect 68600 22512 68900 22568
rect 100 22176 400 22232
rect 68600 21840 68900 21896
rect 100 21504 400 21560
rect 68600 20832 68900 20888
rect 100 20496 400 20552
rect 68600 20160 68900 20216
rect 100 19824 400 19880
rect 68600 19488 68900 19544
rect 100 19152 400 19208
rect 68600 18816 68900 18872
rect 100 18480 400 18536
rect 68600 18144 68900 18200
rect 100 17808 400 17864
rect 68600 17472 68900 17528
rect 100 17136 400 17192
rect 68600 16800 68900 16856
rect 100 16464 400 16520
rect 68600 16128 68900 16184
rect 100 15456 400 15512
rect 68600 15120 68900 15176
rect 100 14784 400 14840
rect 68600 14448 68900 14504
rect 100 14112 400 14168
rect 68600 13776 68900 13832
rect 100 13440 400 13496
rect 68600 13104 68900 13160
rect 100 12768 400 12824
rect 68600 12432 68900 12488
rect 100 12096 400 12152
rect 68600 11760 68900 11816
rect 100 11424 400 11480
rect 68600 11088 68900 11144
rect 100 10752 400 10808
rect 68600 10080 68900 10136
rect 100 9744 400 9800
rect 68600 9408 68900 9464
rect 100 9072 400 9128
rect 68600 8736 68900 8792
rect 100 8400 400 8456
rect 68600 8064 68900 8120
rect 100 7728 400 7784
rect 68600 7392 68900 7448
rect 100 7056 400 7112
rect 68600 6720 68900 6776
rect 100 6384 400 6440
rect 68600 6048 68900 6104
rect 100 5712 400 5768
rect 68600 5376 68900 5432
rect 100 4704 400 4760
rect 68600 4368 68900 4424
rect 100 4032 400 4088
rect 68600 3696 68900 3752
rect 100 3360 400 3416
rect 68600 3024 68900 3080
rect 100 2688 400 2744
rect 68600 2352 68900 2408
rect 100 2016 400 2072
rect 68600 1680 68900 1736
rect 100 1344 400 1400
rect 68600 1008 68900 1064
rect 100 672 400 728
rect 68600 336 68900 392
<< obsm3 >>
rect 9 78374 68978 78414
rect 9 78258 68570 78374
rect 68930 78258 68978 78374
rect 9 78038 68978 78258
rect 9 77922 70 78038
rect 430 77922 68978 78038
rect 9 77702 68978 77922
rect 9 77586 68570 77702
rect 68930 77586 68978 77702
rect 9 77366 68978 77586
rect 9 77250 70 77366
rect 430 77250 68978 77366
rect 9 77030 68978 77250
rect 9 76914 68570 77030
rect 68930 76914 68978 77030
rect 9 76694 68978 76914
rect 9 76578 70 76694
rect 430 76578 68978 76694
rect 9 76358 68978 76578
rect 9 76242 68570 76358
rect 68930 76242 68978 76358
rect 9 76022 68978 76242
rect 9 75906 70 76022
rect 430 75906 68978 76022
rect 9 75686 68978 75906
rect 9 75570 68570 75686
rect 68930 75570 68978 75686
rect 9 75350 68978 75570
rect 9 75234 70 75350
rect 430 75234 68978 75350
rect 9 75014 68978 75234
rect 9 74898 68570 75014
rect 68930 74898 68978 75014
rect 9 74342 68978 74898
rect 9 74226 70 74342
rect 430 74226 68978 74342
rect 9 74006 68978 74226
rect 9 73890 68570 74006
rect 68930 73890 68978 74006
rect 9 73670 68978 73890
rect 9 73554 70 73670
rect 430 73554 68978 73670
rect 9 73334 68978 73554
rect 9 73218 68570 73334
rect 68930 73218 68978 73334
rect 9 72998 68978 73218
rect 9 72882 70 72998
rect 430 72882 68978 72998
rect 9 72662 68978 72882
rect 9 72546 68570 72662
rect 68930 72546 68978 72662
rect 9 72326 68978 72546
rect 9 72210 70 72326
rect 430 72210 68978 72326
rect 9 71990 68978 72210
rect 9 71874 68570 71990
rect 68930 71874 68978 71990
rect 9 71654 68978 71874
rect 9 71538 70 71654
rect 430 71538 68978 71654
rect 9 71318 68978 71538
rect 9 71202 68570 71318
rect 68930 71202 68978 71318
rect 9 70982 68978 71202
rect 9 70866 70 70982
rect 430 70866 68978 70982
rect 9 70646 68978 70866
rect 9 70530 68570 70646
rect 68930 70530 68978 70646
rect 9 70310 68978 70530
rect 9 70194 70 70310
rect 430 70194 68978 70310
rect 9 69974 68978 70194
rect 9 69858 68570 69974
rect 68930 69858 68978 69974
rect 9 69638 68978 69858
rect 9 69522 70 69638
rect 430 69522 68978 69638
rect 9 68966 68978 69522
rect 9 68850 68570 68966
rect 68930 68850 68978 68966
rect 9 68630 68978 68850
rect 9 68514 70 68630
rect 430 68514 68978 68630
rect 9 68294 68978 68514
rect 9 68178 68570 68294
rect 68930 68178 68978 68294
rect 9 67958 68978 68178
rect 9 67842 70 67958
rect 430 67842 68978 67958
rect 9 67622 68978 67842
rect 9 67506 68570 67622
rect 68930 67506 68978 67622
rect 9 67286 68978 67506
rect 9 67170 70 67286
rect 430 67170 68978 67286
rect 9 66950 68978 67170
rect 9 66834 68570 66950
rect 68930 66834 68978 66950
rect 9 66614 68978 66834
rect 9 66498 70 66614
rect 430 66498 68978 66614
rect 9 66278 68978 66498
rect 9 66162 68570 66278
rect 68930 66162 68978 66278
rect 9 65942 68978 66162
rect 9 65826 70 65942
rect 430 65826 68978 65942
rect 9 65606 68978 65826
rect 9 65490 68570 65606
rect 68930 65490 68978 65606
rect 9 65270 68978 65490
rect 9 65154 70 65270
rect 430 65154 68978 65270
rect 9 64934 68978 65154
rect 9 64818 68570 64934
rect 68930 64818 68978 64934
rect 9 64598 68978 64818
rect 9 64482 70 64598
rect 430 64482 68978 64598
rect 9 64262 68978 64482
rect 9 64146 68570 64262
rect 68930 64146 68978 64262
rect 9 63590 68978 64146
rect 9 63474 70 63590
rect 430 63474 68978 63590
rect 9 63254 68978 63474
rect 9 63138 68570 63254
rect 68930 63138 68978 63254
rect 9 62918 68978 63138
rect 9 62802 70 62918
rect 430 62802 68978 62918
rect 9 62582 68978 62802
rect 9 62466 68570 62582
rect 68930 62466 68978 62582
rect 9 62246 68978 62466
rect 9 62130 70 62246
rect 430 62130 68978 62246
rect 9 61910 68978 62130
rect 9 61794 68570 61910
rect 68930 61794 68978 61910
rect 9 61574 68978 61794
rect 9 61458 70 61574
rect 430 61458 68978 61574
rect 9 61238 68978 61458
rect 9 61122 68570 61238
rect 68930 61122 68978 61238
rect 9 60902 68978 61122
rect 9 60786 70 60902
rect 430 60786 68978 60902
rect 9 60566 68978 60786
rect 9 60450 68570 60566
rect 68930 60450 68978 60566
rect 9 60230 68978 60450
rect 9 60114 70 60230
rect 430 60114 68978 60230
rect 9 59894 68978 60114
rect 9 59778 68570 59894
rect 68930 59778 68978 59894
rect 9 59558 68978 59778
rect 9 59442 70 59558
rect 430 59442 68978 59558
rect 9 59222 68978 59442
rect 9 59106 68570 59222
rect 68930 59106 68978 59222
rect 9 58886 68978 59106
rect 9 58770 70 58886
rect 430 58770 68978 58886
rect 9 58214 68978 58770
rect 9 58098 68570 58214
rect 68930 58098 68978 58214
rect 9 57878 68978 58098
rect 9 57762 70 57878
rect 430 57762 68978 57878
rect 9 57542 68978 57762
rect 9 57426 68570 57542
rect 68930 57426 68978 57542
rect 9 57206 68978 57426
rect 9 57090 70 57206
rect 430 57090 68978 57206
rect 9 56870 68978 57090
rect 9 56754 68570 56870
rect 68930 56754 68978 56870
rect 9 56534 68978 56754
rect 9 56418 70 56534
rect 430 56418 68978 56534
rect 9 56198 68978 56418
rect 9 56082 68570 56198
rect 68930 56082 68978 56198
rect 9 55862 68978 56082
rect 9 55746 70 55862
rect 430 55746 68978 55862
rect 9 55526 68978 55746
rect 9 55410 68570 55526
rect 68930 55410 68978 55526
rect 9 55190 68978 55410
rect 9 55074 70 55190
rect 430 55074 68978 55190
rect 9 54854 68978 55074
rect 9 54738 68570 54854
rect 68930 54738 68978 54854
rect 9 54518 68978 54738
rect 9 54402 70 54518
rect 430 54402 68978 54518
rect 9 54182 68978 54402
rect 9 54066 68570 54182
rect 68930 54066 68978 54182
rect 9 53846 68978 54066
rect 9 53730 70 53846
rect 430 53730 68978 53846
rect 9 53510 68978 53730
rect 9 53394 68570 53510
rect 68930 53394 68978 53510
rect 9 52838 68978 53394
rect 9 52722 70 52838
rect 430 52722 68978 52838
rect 9 52502 68978 52722
rect 9 52386 68570 52502
rect 68930 52386 68978 52502
rect 9 52166 68978 52386
rect 9 52050 70 52166
rect 430 52050 68978 52166
rect 9 51830 68978 52050
rect 9 51714 68570 51830
rect 68930 51714 68978 51830
rect 9 51494 68978 51714
rect 9 51378 70 51494
rect 430 51378 68978 51494
rect 9 51158 68978 51378
rect 9 51042 68570 51158
rect 68930 51042 68978 51158
rect 9 50822 68978 51042
rect 9 50706 70 50822
rect 430 50706 68978 50822
rect 9 50486 68978 50706
rect 9 50370 68570 50486
rect 68930 50370 68978 50486
rect 9 50150 68978 50370
rect 9 50034 70 50150
rect 430 50034 68978 50150
rect 9 49814 68978 50034
rect 9 49698 68570 49814
rect 68930 49698 68978 49814
rect 9 49478 68978 49698
rect 9 49362 70 49478
rect 430 49362 68978 49478
rect 9 49142 68978 49362
rect 9 49026 68570 49142
rect 68930 49026 68978 49142
rect 9 48806 68978 49026
rect 9 48690 70 48806
rect 430 48690 68978 48806
rect 9 48470 68978 48690
rect 9 48354 68570 48470
rect 68930 48354 68978 48470
rect 9 48134 68978 48354
rect 9 48018 70 48134
rect 430 48018 68978 48134
rect 9 47462 68978 48018
rect 9 47346 68570 47462
rect 68930 47346 68978 47462
rect 9 47126 68978 47346
rect 9 47010 70 47126
rect 430 47010 68978 47126
rect 9 46790 68978 47010
rect 9 46674 68570 46790
rect 68930 46674 68978 46790
rect 9 46454 68978 46674
rect 9 46338 70 46454
rect 430 46338 68978 46454
rect 9 46118 68978 46338
rect 9 46002 68570 46118
rect 68930 46002 68978 46118
rect 9 45782 68978 46002
rect 9 45666 70 45782
rect 430 45666 68978 45782
rect 9 45446 68978 45666
rect 9 45330 68570 45446
rect 68930 45330 68978 45446
rect 9 45110 68978 45330
rect 9 44994 70 45110
rect 430 44994 68978 45110
rect 9 44774 68978 44994
rect 9 44658 68570 44774
rect 68930 44658 68978 44774
rect 9 44438 68978 44658
rect 9 44322 70 44438
rect 430 44322 68978 44438
rect 9 44102 68978 44322
rect 9 43986 68570 44102
rect 68930 43986 68978 44102
rect 9 43766 68978 43986
rect 9 43650 70 43766
rect 430 43650 68978 43766
rect 9 43430 68978 43650
rect 9 43314 68570 43430
rect 68930 43314 68978 43430
rect 9 43094 68978 43314
rect 9 42978 70 43094
rect 430 42978 68978 43094
rect 9 42758 68978 42978
rect 9 42642 68570 42758
rect 68930 42642 68978 42758
rect 9 42086 68978 42642
rect 9 41970 70 42086
rect 430 41970 68978 42086
rect 9 41750 68978 41970
rect 9 41634 68570 41750
rect 68930 41634 68978 41750
rect 9 41414 68978 41634
rect 9 41298 70 41414
rect 430 41298 68978 41414
rect 9 41078 68978 41298
rect 9 40962 68570 41078
rect 68930 40962 68978 41078
rect 9 40742 68978 40962
rect 9 40626 70 40742
rect 430 40626 68978 40742
rect 9 40406 68978 40626
rect 9 40290 68570 40406
rect 68930 40290 68978 40406
rect 9 40070 68978 40290
rect 9 39954 70 40070
rect 430 39954 68978 40070
rect 9 39734 68978 39954
rect 9 39618 68570 39734
rect 68930 39618 68978 39734
rect 9 39398 68978 39618
rect 9 39282 70 39398
rect 430 39282 68978 39398
rect 9 39062 68978 39282
rect 9 38946 68570 39062
rect 68930 38946 68978 39062
rect 9 38726 68978 38946
rect 9 38610 70 38726
rect 430 38610 68978 38726
rect 9 38390 68978 38610
rect 9 38274 68570 38390
rect 68930 38274 68978 38390
rect 9 38054 68978 38274
rect 9 37938 70 38054
rect 430 37938 68978 38054
rect 9 37718 68978 37938
rect 9 37602 68570 37718
rect 68930 37602 68978 37718
rect 9 37046 68978 37602
rect 9 36930 70 37046
rect 430 36930 68978 37046
rect 9 36710 68978 36930
rect 9 36594 68570 36710
rect 68930 36594 68978 36710
rect 9 36374 68978 36594
rect 9 36258 70 36374
rect 430 36258 68978 36374
rect 9 36038 68978 36258
rect 9 35922 68570 36038
rect 68930 35922 68978 36038
rect 9 35702 68978 35922
rect 9 35586 70 35702
rect 430 35586 68978 35702
rect 9 35366 68978 35586
rect 9 35250 68570 35366
rect 68930 35250 68978 35366
rect 9 35030 68978 35250
rect 9 34914 70 35030
rect 430 34914 68978 35030
rect 9 34694 68978 34914
rect 9 34578 68570 34694
rect 68930 34578 68978 34694
rect 9 34358 68978 34578
rect 9 34242 70 34358
rect 430 34242 68978 34358
rect 9 34022 68978 34242
rect 9 33906 68570 34022
rect 68930 33906 68978 34022
rect 9 33686 68978 33906
rect 9 33570 70 33686
rect 430 33570 68978 33686
rect 9 33350 68978 33570
rect 9 33234 68570 33350
rect 68930 33234 68978 33350
rect 9 33014 68978 33234
rect 9 32898 70 33014
rect 430 32898 68978 33014
rect 9 32678 68978 32898
rect 9 32562 68570 32678
rect 68930 32562 68978 32678
rect 9 32342 68978 32562
rect 9 32226 70 32342
rect 430 32226 68978 32342
rect 9 31670 68978 32226
rect 9 31554 68570 31670
rect 68930 31554 68978 31670
rect 9 31334 68978 31554
rect 9 31218 70 31334
rect 430 31218 68978 31334
rect 9 30998 68978 31218
rect 9 30882 68570 30998
rect 68930 30882 68978 30998
rect 9 30662 68978 30882
rect 9 30546 70 30662
rect 430 30546 68978 30662
rect 9 30326 68978 30546
rect 9 30210 68570 30326
rect 68930 30210 68978 30326
rect 9 29990 68978 30210
rect 9 29874 70 29990
rect 430 29874 68978 29990
rect 9 29654 68978 29874
rect 9 29538 68570 29654
rect 68930 29538 68978 29654
rect 9 29318 68978 29538
rect 9 29202 70 29318
rect 430 29202 68978 29318
rect 9 28982 68978 29202
rect 9 28866 68570 28982
rect 68930 28866 68978 28982
rect 9 28646 68978 28866
rect 9 28530 70 28646
rect 430 28530 68978 28646
rect 9 28310 68978 28530
rect 9 28194 68570 28310
rect 68930 28194 68978 28310
rect 9 27974 68978 28194
rect 9 27858 70 27974
rect 430 27858 68978 27974
rect 9 27638 68978 27858
rect 9 27522 68570 27638
rect 68930 27522 68978 27638
rect 9 27302 68978 27522
rect 9 27186 70 27302
rect 430 27186 68978 27302
rect 9 26966 68978 27186
rect 9 26850 68570 26966
rect 68930 26850 68978 26966
rect 9 26294 68978 26850
rect 9 26178 70 26294
rect 430 26178 68978 26294
rect 9 25958 68978 26178
rect 9 25842 68570 25958
rect 68930 25842 68978 25958
rect 9 25622 68978 25842
rect 9 25506 70 25622
rect 430 25506 68978 25622
rect 9 25286 68978 25506
rect 9 25170 68570 25286
rect 68930 25170 68978 25286
rect 9 24950 68978 25170
rect 9 24834 70 24950
rect 430 24834 68978 24950
rect 9 24614 68978 24834
rect 9 24498 68570 24614
rect 68930 24498 68978 24614
rect 9 24278 68978 24498
rect 9 24162 70 24278
rect 430 24162 68978 24278
rect 9 23942 68978 24162
rect 9 23826 68570 23942
rect 68930 23826 68978 23942
rect 9 23606 68978 23826
rect 9 23490 70 23606
rect 430 23490 68978 23606
rect 9 23270 68978 23490
rect 9 23154 68570 23270
rect 68930 23154 68978 23270
rect 9 22934 68978 23154
rect 9 22818 70 22934
rect 430 22818 68978 22934
rect 9 22598 68978 22818
rect 9 22482 68570 22598
rect 68930 22482 68978 22598
rect 9 22262 68978 22482
rect 9 22146 70 22262
rect 430 22146 68978 22262
rect 9 21926 68978 22146
rect 9 21810 68570 21926
rect 68930 21810 68978 21926
rect 9 21590 68978 21810
rect 9 21474 70 21590
rect 430 21474 68978 21590
rect 9 20918 68978 21474
rect 9 20802 68570 20918
rect 68930 20802 68978 20918
rect 9 20582 68978 20802
rect 9 20466 70 20582
rect 430 20466 68978 20582
rect 9 20246 68978 20466
rect 9 20130 68570 20246
rect 68930 20130 68978 20246
rect 9 19910 68978 20130
rect 9 19794 70 19910
rect 430 19794 68978 19910
rect 9 19574 68978 19794
rect 9 19458 68570 19574
rect 68930 19458 68978 19574
rect 9 19238 68978 19458
rect 9 19122 70 19238
rect 430 19122 68978 19238
rect 9 18902 68978 19122
rect 9 18786 68570 18902
rect 68930 18786 68978 18902
rect 9 18566 68978 18786
rect 9 18450 70 18566
rect 430 18450 68978 18566
rect 9 18230 68978 18450
rect 9 18114 68570 18230
rect 68930 18114 68978 18230
rect 9 17894 68978 18114
rect 9 17778 70 17894
rect 430 17778 68978 17894
rect 9 17558 68978 17778
rect 9 17442 68570 17558
rect 68930 17442 68978 17558
rect 9 17222 68978 17442
rect 9 17106 70 17222
rect 430 17106 68978 17222
rect 9 16886 68978 17106
rect 9 16770 68570 16886
rect 68930 16770 68978 16886
rect 9 16550 68978 16770
rect 9 16434 70 16550
rect 430 16434 68978 16550
rect 9 16214 68978 16434
rect 9 16098 68570 16214
rect 68930 16098 68978 16214
rect 9 15542 68978 16098
rect 9 15426 70 15542
rect 430 15426 68978 15542
rect 9 15206 68978 15426
rect 9 15090 68570 15206
rect 68930 15090 68978 15206
rect 9 14870 68978 15090
rect 9 14754 70 14870
rect 430 14754 68978 14870
rect 9 14534 68978 14754
rect 9 14418 68570 14534
rect 68930 14418 68978 14534
rect 9 14198 68978 14418
rect 9 14082 70 14198
rect 430 14082 68978 14198
rect 9 13862 68978 14082
rect 9 13746 68570 13862
rect 68930 13746 68978 13862
rect 9 13526 68978 13746
rect 9 13410 70 13526
rect 430 13410 68978 13526
rect 9 13190 68978 13410
rect 9 13074 68570 13190
rect 68930 13074 68978 13190
rect 9 12854 68978 13074
rect 9 12738 70 12854
rect 430 12738 68978 12854
rect 9 12518 68978 12738
rect 9 12402 68570 12518
rect 68930 12402 68978 12518
rect 9 12182 68978 12402
rect 9 12066 70 12182
rect 430 12066 68978 12182
rect 9 11846 68978 12066
rect 9 11730 68570 11846
rect 68930 11730 68978 11846
rect 9 11510 68978 11730
rect 9 11394 70 11510
rect 430 11394 68978 11510
rect 9 11174 68978 11394
rect 9 11058 68570 11174
rect 68930 11058 68978 11174
rect 9 10838 68978 11058
rect 9 10722 70 10838
rect 430 10722 68978 10838
rect 9 10166 68978 10722
rect 9 10050 68570 10166
rect 68930 10050 68978 10166
rect 9 9830 68978 10050
rect 9 9714 70 9830
rect 430 9714 68978 9830
rect 9 9494 68978 9714
rect 9 9378 68570 9494
rect 68930 9378 68978 9494
rect 9 9158 68978 9378
rect 9 9042 70 9158
rect 430 9042 68978 9158
rect 9 8822 68978 9042
rect 9 8706 68570 8822
rect 68930 8706 68978 8822
rect 9 8486 68978 8706
rect 9 8370 70 8486
rect 430 8370 68978 8486
rect 9 8150 68978 8370
rect 9 8034 68570 8150
rect 68930 8034 68978 8150
rect 9 7814 68978 8034
rect 9 7698 70 7814
rect 430 7698 68978 7814
rect 9 7478 68978 7698
rect 9 7362 68570 7478
rect 68930 7362 68978 7478
rect 9 7142 68978 7362
rect 9 7026 70 7142
rect 430 7026 68978 7142
rect 9 6806 68978 7026
rect 9 6690 68570 6806
rect 68930 6690 68978 6806
rect 9 6470 68978 6690
rect 9 6354 70 6470
rect 430 6354 68978 6470
rect 9 6134 68978 6354
rect 9 6018 68570 6134
rect 68930 6018 68978 6134
rect 9 5798 68978 6018
rect 9 5682 70 5798
rect 430 5682 68978 5798
rect 9 5462 68978 5682
rect 9 5346 68570 5462
rect 68930 5346 68978 5462
rect 9 4790 68978 5346
rect 9 4674 70 4790
rect 430 4674 68978 4790
rect 9 4454 68978 4674
rect 9 4338 68570 4454
rect 68930 4338 68978 4454
rect 9 4118 68978 4338
rect 9 4002 70 4118
rect 430 4002 68978 4118
rect 9 3782 68978 4002
rect 9 3666 68570 3782
rect 68930 3666 68978 3782
rect 9 3446 68978 3666
rect 9 3330 70 3446
rect 430 3330 68978 3446
rect 9 3110 68978 3330
rect 9 2994 68570 3110
rect 68930 2994 68978 3110
rect 9 2774 68978 2994
rect 9 2658 70 2774
rect 430 2658 68978 2774
rect 9 2438 68978 2658
rect 9 2322 68570 2438
rect 68930 2322 68978 2438
rect 9 2102 68978 2322
rect 9 1986 70 2102
rect 430 1986 68978 2102
rect 9 1766 68978 1986
rect 9 1650 68570 1766
rect 68930 1650 68978 1766
rect 9 1430 68978 1650
rect 9 1314 70 1430
rect 430 1314 68978 1430
rect 9 1094 68978 1314
rect 9 978 68570 1094
rect 68930 978 68978 1094
rect 9 758 68978 978
rect 9 642 70 758
rect 430 642 68978 758
rect 9 422 68978 642
rect 9 350 68570 422
rect 68930 350 68978 422
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
<< obsm4 >>
rect 1862 1508 2194 76543
rect 2414 1508 9874 76543
rect 10094 1508 17554 76543
rect 17774 1508 25234 76543
rect 25454 1508 32914 76543
rect 33134 1508 40594 76543
rect 40814 1508 48274 76543
rect 48494 1508 55954 76543
rect 56174 1508 63634 76543
rect 63854 1508 66178 76543
rect 1862 1353 66178 1508
<< labels >>
rlabel metal3 s 100 51408 400 51464 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 52080 400 52136 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 25536 400 25592 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 45024 400 45080 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 30576 400 30632 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 26208 400 26264 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 33936 79600 33992 79900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 68600 20160 68900 20216 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 68600 75600 68900 75656 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 44688 79600 44744 79900 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 68600 3696 68900 3752 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3696 79600 3752 79900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 54096 79600 54152 79900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 52080 100 52136 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 68880 79600 68936 79900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 68600 69888 68900 69944 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 61488 100 61544 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 62160 400 62216 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 50736 400 50792 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 57792 400 57848 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 46368 400 46424 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 68600 78960 68900 79016 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 48720 100 48776 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 31248 400 31304 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 62832 100 62888 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 7728 400 7784 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 100 66528 400 66584 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 61152 79600 61208 79900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 68600 71232 68900 71288 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 68600 61824 68900 61880 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 68600 78288 68900 78344 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 68600 38976 68900 39032 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 14112 400 14168 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 68600 19488 68900 19544 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 55440 79600 55496 79900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 34272 400 34328 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 38640 400 38696 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 68600 57456 68900 57512 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 68600 53424 68900 53480 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 100 77280 400 77336 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 45696 100 45752 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 19152 400 19208 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 67872 100 67928 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 41664 79600 41720 79900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 21504 100 21560 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 7056 100 7112 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 77952 400 78008 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 20832 79600 20888 79900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 14448 79600 14504 79900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 37632 79600 37688 79900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 63504 100 63560 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 68600 24528 68900 24584 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 66864 79600 66920 79900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 21504 400 21560 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 10752 400 10808 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 100 67872 400 67928 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 62160 100 62216 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 100 75936 400 75992 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 68600 43344 68900 43400 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 68600 33936 68900 33992 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 68600 1008 68900 1064 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 22848 400 22904 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 59808 79600 59864 79900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 68600 17472 68900 17528 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 60816 400 60872 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 68600 72576 68900 72632 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 35952 79600 36008 79900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 68600 35280 68900 35336 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 55776 400 55832 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 9744 400 9800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 49056 79600 49112 79900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 58800 400 58856 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 30240 79600 30296 79900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 36960 400 37016 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 68600 77616 68900 77672 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6720 79600 6776 79900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 17472 79600 17528 79900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 48048 100 48104 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 67536 79600 67592 79900 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 74256 400 74312 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 55104 400 55160 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 29904 100 29960 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 68600 67536 68900 67592 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 8400 100 8456 400 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 68600 336 68900 392 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 11088 79600 11144 79900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4704 100 4760 400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 68600 12432 68900 12488 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 49392 400 49448 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 68600 21840 68900 21896 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 27888 400 27944 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 65184 100 65240 400 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 68600 7392 68900 7448 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 31248 100 31304 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 24864 100 24920 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 46704 79600 46760 79900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 50736 100 50792 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 68600 31584 68900 31640 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 62496 79600 62552 79900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 26208 100 26264 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 40992 79600 41048 79900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 27216 400 27272 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 49392 100 49448 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 44352 100 44408 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 17808 100 17864 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 3360 400 3416 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 28896 79600 28952 79900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 34272 100 34328 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 25872 79600 25928 79900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 13440 400 13496 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 42000 400 42056 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 54432 100 54488 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 19152 100 19208 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 37968 400 38024 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 68600 74928 68900 74984 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 68600 38304 68900 38360 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 22848 100 22904 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 24528 79600 24584 79900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 100 65184 400 65240 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 68600 59136 68900 59192 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 1680 79600 1736 79900 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 68600 16800 68900 16856 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 31584 79600 31640 79900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 11424 400 11480 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 11760 79600 11816 79900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 68600 20832 68900 20888 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 56448 400 56504 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 32928 400 32984 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 68600 61152 68900 61208 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 32592 79600 32648 79900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 10080 79600 10136 79900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 40320 79600 40376 79900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 100 67200 400 67256 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 70224 400 70280 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 68600 23856 68900 23912 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 27552 79600 27608 79900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 5712 400 5768 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 57456 79600 57512 79900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 29904 400 29960 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 50064 400 50120 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 336 79600 392 79900 6 la_data_in[34]
port 142 nsew signal input
rlabel metal3 s 100 65856 400 65912 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 52752 100 52808 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal3 s 100 72912 400 72968 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 33600 100 33656 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 35280 79600 35336 79900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 68600 46032 68900 46088 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 25536 100 25592 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 35616 100 35672 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 64848 79600 64904 79900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 68600 6048 68900 6104 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 24192 100 24248 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 68600 59808 68900 59864 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 46368 100 46424 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 29568 79600 29624 79900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 23184 79600 23240 79900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 1008 79600 1064 79900 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 23856 79600 23912 79900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 34944 100 35000 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 68600 30240 68900 30296 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 52416 79600 52472 79900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 47376 79600 47432 79900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 19824 400 19880 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 22176 400 22232 6 la_data_in[56]
port 166 nsew signal input
rlabel metal3 s 100 76608 400 76664 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 27216 100 27272 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 68600 73248 68900 73304 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 12768 100 12824 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 68600 54768 68900 54824 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 2016 400 2072 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 43680 100 43736 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 13776 79600 13832 79900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 14784 100 14840 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 68600 32592 68900 32648 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1344 400 1400 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 61824 79600 61880 79900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 59136 79600 59192 79900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 68600 45360 68900 45416 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 53760 400 53816 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 27888 100 27944 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 68600 35952 68900 36008 6 la_data_out[14]
port 184 nsew signal output
rlabel metal3 s 100 63504 400 63560 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 68600 46704 68900 46760 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 30912 79600 30968 79900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 68600 66864 68900 66920 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 39312 100 39368 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 68600 40320 68900 40376 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 68600 16128 68900 16184 6 la_data_out[20]
port 191 nsew signal output
rlabel metal3 s 100 73584 400 73640 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 68600 51744 68900 51800 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 22176 100 22232 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 33600 400 33656 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 39984 100 40040 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 72240 400 72296 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 39648 79600 39704 79900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 68600 64848 68900 64904 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 32256 100 32312 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 17136 400 17192 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 68600 39648 68900 39704 6 la_data_out[30]
port 202 nsew signal output
rlabel metal3 s 68600 8736 68900 8792 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 38304 79600 38360 79900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 68600 18816 68900 18872 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 36288 100 36344 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 34608 79600 34664 79900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 68600 65520 68900 65576 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 68600 34608 68900 34664 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 68600 6720 68900 6776 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 68600 15120 68900 15176 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 12096 400 12152 6 la_data_out[3]
port 212 nsew signal output
rlabel metal3 s 68600 3024 68900 3080 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 68600 28224 68900 28280 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 68600 68208 68900 68264 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 4032 100 4088 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 30576 100 30632 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 6048 79600 6104 79900 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 5376 79600 5432 79900 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 52752 400 52808 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 17136 100 17192 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 67200 100 67256 400 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 36624 79600 36680 79900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 20160 79600 20216 79900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal3 s 100 71568 400 71624 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 68600 10080 68900 10136 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 70896 400 70952 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 68600 56112 68900 56168 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 22512 79600 22568 79900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 68600 23184 68900 23240 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 51072 79600 51128 79900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 68600 56784 68900 56840 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 28560 400 28616 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 68600 49728 68900 49784 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 54768 79600 54824 79900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 19824 100 19880 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 64512 100 64568 400 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 68600 11088 68900 11144 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 68600 26880 68900 26936 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 66192 79600 66248 79900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 4032 400 4088 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 68600 40992 68900 41048 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 68600 33264 68900 33320 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 68600 58128 68900 58184 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 68600 47376 68900 47432 6 la_oenb[11]
port 245 nsew signal input
rlabel metal3 s 100 75264 400 75320 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 59472 400 59528 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 55104 100 55160 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 65856 100 65912 400 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 10752 100 10808 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 9072 400 9128 6 la_oenb[17]
port 251 nsew signal input
rlabel metal3 s 100 79296 400 79352 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 68600 11760 68900 11816 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 8736 79600 8792 79900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 25200 79600 25256 79900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 49728 79600 49784 79900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 20496 100 20552 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 68600 51072 68900 51128 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 66528 100 66584 400 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 9408 79600 9464 79900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 13440 100 13496 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 45696 400 45752 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 68600 76272 68900 76328 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 68208 79600 68264 79900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 68600 68880 68900 68936 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 26880 79600 26936 79900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 68600 66192 68900 66248 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 37968 100 38024 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 7392 79600 7448 79900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 2016 100 2072 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 672 100 728 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 4368 79600 4424 79900 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 38640 100 38696 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 32256 400 32312 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 40656 400 40712 6 la_oenb[3]
port 276 nsew signal input
rlabel metal3 s 68600 14448 68900 14504 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 21840 79600 21896 79900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 47040 400 47096 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 14112 100 14168 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 32928 100 32984 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 56112 79600 56168 79900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 59472 100 59528 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 8400 400 8456 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 672 400 728 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 100 69552 400 69608 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 57120 100 57176 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 18816 79600 18872 79900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal3 s 68600 4368 68900 4424 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 68600 52416 68900 52472 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 39984 400 40040 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 68600 44016 68900 44072 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 56448 100 56504 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 60480 79600 60536 79900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal3 s 68600 13104 68900 13160 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 38976 79600 39032 79900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 68544 100 68600 400 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 36288 400 36344 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 9072 100 9128 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 68600 42672 68900 42728 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 17808 400 17864 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 68600 54096 68900 54152 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 18480 100 18536 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal3 s 68600 1680 68900 1736 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 16128 79600 16184 79900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 58128 79600 58184 79900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 68600 62496 68900 62552 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 13104 79600 13160 79900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 48048 400 48104 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 68600 18144 68900 18200 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 8064 79600 8120 79900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 68600 30912 68900 30968 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 44016 79600 44072 79900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 28224 79600 28280 79900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 43008 400 43064 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 6384 100 6440 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 41328 100 41384 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 7056 400 7112 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 68600 55440 68900 55496 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 47040 100 47096 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 41328 400 41384 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 68600 28896 68900 28952 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 68600 2352 68900 2408 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 4704 400 4760 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 64176 79600 64232 79900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 42000 100 42056 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 60144 100 60200 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 68600 22512 68900 22568 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 3024 79600 3080 79900 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 12768 400 12824 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 7728 100 7784 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 19488 79600 19544 79900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 68600 49056 68900 49112 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 68600 76944 68900 77000 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 29232 100 29288 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 29232 400 29288 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 68600 36624 68900 36680 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 57792 100 57848 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 51744 79600 51800 79900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 55776 100 55832 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 18480 400 18536 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 3360 100 3416 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal3 s 68600 5376 68900 5432 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 68600 25200 68900 25256 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 18144 79600 18200 79900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 68600 70560 68900 70616 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 57120 400 57176 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal3 s 100 62832 400 62888 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 60144 400 60200 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 15456 400 15512 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 68600 44688 68900 44744 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 43008 100 43064 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 45360 79600 45416 79900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 63168 79600 63224 79900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal3 s 100 78624 400 78680 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 11424 100 11480 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 34944 400 35000 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 65520 79600 65576 79900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 44352 400 44408 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 68600 64176 68900 64232 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 68600 29568 68900 29624 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 51408 100 51464 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 56784 79600 56840 79900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 12432 79600 12488 79900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 23520 100 23576 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 68600 50400 68900 50456 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 60816 100 60872 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 68600 27552 68900 27608 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal3 s 68600 8064 68900 8120 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 12096 100 12152 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 37296 100 37352 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 68600 37632 68900 37688 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 53424 79600 53480 79900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 68600 71904 68900 71960 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal3 s 68600 9408 68900 9464 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 14784 400 14840 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 68600 48384 68900 48440 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1344 100 1400 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 68600 73920 68900 73976 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 50400 79600 50456 79900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal3 s 68600 13776 68900 13832 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 48384 79600 48440 79900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 20496 400 20552 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 23520 400 23576 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 50064 100 50120 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 58800 100 58856 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 35616 400 35672 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal3 s 100 64512 400 64568 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 15120 79600 15176 79900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 24192 400 24248 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 15456 100 15512 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 5712 100 5768 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 33264 79600 33320 79900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 16800 79600 16856 79900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 40656 100 40712 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 46032 79600 46088 79900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 68600 25872 68900 25928 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 48720 400 48776 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 68600 63168 68900 63224 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 16464 100 16520 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 28560 100 28616 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 6384 400 6440 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 68600 60480 68900 60536 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 45024 100 45080 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 43344 79600 43400 79900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 42672 79600 42728 79900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal3 s 100 68544 400 68600 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 2352 79600 2408 79900 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 53760 100 53816 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 16464 400 16520 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 61488 400 61544 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 68600 41664 68900 41720 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 69000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18720374
string GDS_FILE /home/runner/work/gf180-mpw0-serv/gf180-mpw0-serv/openlane/tiny_user_project/runs/22_12_03_00_36/results/signoff/tiny_user_project.magic.gds
string GDS_START 297750
<< end >>

