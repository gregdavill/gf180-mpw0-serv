magic
tech gf180mcuC
magscale 1 5
timestamp 1669991585
<< obsm1 >>
rect 672 855 77663 106329
<< metal2 >>
rect 0 107600 56 107900
rect 672 107600 728 107900
rect 1680 107600 1736 107900
rect 2688 107600 2744 107900
rect 3360 107600 3416 107900
rect 4368 107600 4424 107900
rect 5376 107600 5432 107900
rect 6048 107600 6104 107900
rect 7056 107600 7112 107900
rect 8064 107600 8120 107900
rect 8736 107600 8792 107900
rect 9744 107600 9800 107900
rect 10752 107600 10808 107900
rect 11424 107600 11480 107900
rect 12432 107600 12488 107900
rect 13440 107600 13496 107900
rect 14112 107600 14168 107900
rect 15120 107600 15176 107900
rect 16128 107600 16184 107900
rect 16800 107600 16856 107900
rect 17808 107600 17864 107900
rect 18816 107600 18872 107900
rect 19488 107600 19544 107900
rect 20496 107600 20552 107900
rect 21504 107600 21560 107900
rect 22176 107600 22232 107900
rect 23184 107600 23240 107900
rect 24192 107600 24248 107900
rect 24864 107600 24920 107900
rect 25872 107600 25928 107900
rect 26880 107600 26936 107900
rect 27552 107600 27608 107900
rect 28560 107600 28616 107900
rect 29568 107600 29624 107900
rect 30240 107600 30296 107900
rect 31248 107600 31304 107900
rect 32256 107600 32312 107900
rect 32928 107600 32984 107900
rect 33936 107600 33992 107900
rect 34944 107600 35000 107900
rect 35616 107600 35672 107900
rect 36624 107600 36680 107900
rect 37632 107600 37688 107900
rect 38304 107600 38360 107900
rect 39312 107600 39368 107900
rect 40320 107600 40376 107900
rect 40992 107600 41048 107900
rect 42000 107600 42056 107900
rect 43008 107600 43064 107900
rect 43680 107600 43736 107900
rect 44688 107600 44744 107900
rect 45696 107600 45752 107900
rect 46368 107600 46424 107900
rect 47376 107600 47432 107900
rect 48384 107600 48440 107900
rect 49056 107600 49112 107900
rect 50064 107600 50120 107900
rect 51072 107600 51128 107900
rect 51744 107600 51800 107900
rect 52752 107600 52808 107900
rect 53760 107600 53816 107900
rect 54432 107600 54488 107900
rect 55440 107600 55496 107900
rect 56448 107600 56504 107900
rect 57120 107600 57176 107900
rect 58128 107600 58184 107900
rect 59136 107600 59192 107900
rect 59808 107600 59864 107900
rect 60816 107600 60872 107900
rect 61824 107600 61880 107900
rect 62496 107600 62552 107900
rect 63504 107600 63560 107900
rect 64512 107600 64568 107900
rect 65184 107600 65240 107900
rect 66192 107600 66248 107900
rect 67200 107600 67256 107900
rect 67872 107600 67928 107900
rect 68880 107600 68936 107900
rect 69888 107600 69944 107900
rect 70560 107600 70616 107900
rect 71568 107600 71624 107900
rect 72576 107600 72632 107900
rect 73248 107600 73304 107900
rect 74256 107600 74312 107900
rect 75264 107600 75320 107900
rect 75936 107600 75992 107900
rect 76944 107600 77000 107900
rect 77616 107600 77672 107900
rect 0 100 56 400
rect 672 100 728 400
rect 1680 100 1736 400
rect 2352 100 2408 400
rect 3360 100 3416 400
rect 4368 100 4424 400
rect 5040 100 5096 400
rect 6048 100 6104 400
rect 7056 100 7112 400
rect 7728 100 7784 400
rect 8736 100 8792 400
rect 9744 100 9800 400
rect 10416 100 10472 400
rect 11424 100 11480 400
rect 12432 100 12488 400
rect 13104 100 13160 400
rect 14112 100 14168 400
rect 15120 100 15176 400
rect 15792 100 15848 400
rect 16800 100 16856 400
rect 17808 100 17864 400
rect 18480 100 18536 400
rect 19488 100 19544 400
rect 20496 100 20552 400
rect 21168 100 21224 400
rect 22176 100 22232 400
rect 23184 100 23240 400
rect 23856 100 23912 400
rect 24864 100 24920 400
rect 25872 100 25928 400
rect 26544 100 26600 400
rect 27552 100 27608 400
rect 28560 100 28616 400
rect 29232 100 29288 400
rect 30240 100 30296 400
rect 31248 100 31304 400
rect 31920 100 31976 400
rect 32928 100 32984 400
rect 33936 100 33992 400
rect 34608 100 34664 400
rect 35616 100 35672 400
rect 36624 100 36680 400
rect 37296 100 37352 400
rect 38304 100 38360 400
rect 39312 100 39368 400
rect 39984 100 40040 400
rect 40992 100 41048 400
rect 42000 100 42056 400
rect 42672 100 42728 400
rect 43680 100 43736 400
rect 44688 100 44744 400
rect 45360 100 45416 400
rect 46368 100 46424 400
rect 47376 100 47432 400
rect 48048 100 48104 400
rect 49056 100 49112 400
rect 50064 100 50120 400
rect 50736 100 50792 400
rect 51744 100 51800 400
rect 52752 100 52808 400
rect 53424 100 53480 400
rect 54432 100 54488 400
rect 55440 100 55496 400
rect 56112 100 56168 400
rect 57120 100 57176 400
rect 58128 100 58184 400
rect 58800 100 58856 400
rect 59808 100 59864 400
rect 60816 100 60872 400
rect 61488 100 61544 400
rect 62496 100 62552 400
rect 63504 100 63560 400
rect 64176 100 64232 400
rect 65184 100 65240 400
rect 66192 100 66248 400
rect 66864 100 66920 400
rect 67872 100 67928 400
rect 68880 100 68936 400
rect 69552 100 69608 400
rect 70560 100 70616 400
rect 71568 100 71624 400
rect 72240 100 72296 400
rect 73248 100 73304 400
rect 74256 100 74312 400
rect 74928 100 74984 400
rect 75936 100 75992 400
rect 76944 100 77000 400
rect 77616 100 77672 400
<< obsm2 >>
rect 86 107570 642 107600
rect 758 107570 1650 107600
rect 1766 107570 2658 107600
rect 2774 107570 3330 107600
rect 3446 107570 4338 107600
rect 4454 107570 5346 107600
rect 5462 107570 6018 107600
rect 6134 107570 7026 107600
rect 7142 107570 8034 107600
rect 8150 107570 8706 107600
rect 8822 107570 9714 107600
rect 9830 107570 10722 107600
rect 10838 107570 11394 107600
rect 11510 107570 12402 107600
rect 12518 107570 13410 107600
rect 13526 107570 14082 107600
rect 14198 107570 15090 107600
rect 15206 107570 16098 107600
rect 16214 107570 16770 107600
rect 16886 107570 17778 107600
rect 17894 107570 18786 107600
rect 18902 107570 19458 107600
rect 19574 107570 20466 107600
rect 20582 107570 21474 107600
rect 21590 107570 22146 107600
rect 22262 107570 23154 107600
rect 23270 107570 24162 107600
rect 24278 107570 24834 107600
rect 24950 107570 25842 107600
rect 25958 107570 26850 107600
rect 26966 107570 27522 107600
rect 27638 107570 28530 107600
rect 28646 107570 29538 107600
rect 29654 107570 30210 107600
rect 30326 107570 31218 107600
rect 31334 107570 32226 107600
rect 32342 107570 32898 107600
rect 33014 107570 33906 107600
rect 34022 107570 34914 107600
rect 35030 107570 35586 107600
rect 35702 107570 36594 107600
rect 36710 107570 37602 107600
rect 37718 107570 38274 107600
rect 38390 107570 39282 107600
rect 39398 107570 40290 107600
rect 40406 107570 40962 107600
rect 41078 107570 41970 107600
rect 42086 107570 42978 107600
rect 43094 107570 43650 107600
rect 43766 107570 44658 107600
rect 44774 107570 45666 107600
rect 45782 107570 46338 107600
rect 46454 107570 47346 107600
rect 47462 107570 48354 107600
rect 48470 107570 49026 107600
rect 49142 107570 50034 107600
rect 50150 107570 51042 107600
rect 51158 107570 51714 107600
rect 51830 107570 52722 107600
rect 52838 107570 53730 107600
rect 53846 107570 54402 107600
rect 54518 107570 55410 107600
rect 55526 107570 56418 107600
rect 56534 107570 57090 107600
rect 57206 107570 58098 107600
rect 58214 107570 59106 107600
rect 59222 107570 59778 107600
rect 59894 107570 60786 107600
rect 60902 107570 61794 107600
rect 61910 107570 62466 107600
rect 62582 107570 63474 107600
rect 63590 107570 64482 107600
rect 64598 107570 65154 107600
rect 65270 107570 66162 107600
rect 66278 107570 67170 107600
rect 67286 107570 67842 107600
rect 67958 107570 68850 107600
rect 68966 107570 69858 107600
rect 69974 107570 70530 107600
rect 70646 107570 71538 107600
rect 71654 107570 72546 107600
rect 72662 107570 73218 107600
rect 73334 107570 74226 107600
rect 74342 107570 75234 107600
rect 75350 107570 75906 107600
rect 76022 107570 76914 107600
rect 77030 107570 77586 107600
rect 14 430 77658 107570
rect 86 400 642 430
rect 758 400 1650 430
rect 1766 400 2322 430
rect 2438 400 3330 430
rect 3446 400 4338 430
rect 4454 400 5010 430
rect 5126 400 6018 430
rect 6134 400 7026 430
rect 7142 400 7698 430
rect 7814 400 8706 430
rect 8822 400 9714 430
rect 9830 400 10386 430
rect 10502 400 11394 430
rect 11510 400 12402 430
rect 12518 400 13074 430
rect 13190 400 14082 430
rect 14198 400 15090 430
rect 15206 400 15762 430
rect 15878 400 16770 430
rect 16886 400 17778 430
rect 17894 400 18450 430
rect 18566 400 19458 430
rect 19574 400 20466 430
rect 20582 400 21138 430
rect 21254 400 22146 430
rect 22262 400 23154 430
rect 23270 400 23826 430
rect 23942 400 24834 430
rect 24950 400 25842 430
rect 25958 400 26514 430
rect 26630 400 27522 430
rect 27638 400 28530 430
rect 28646 400 29202 430
rect 29318 400 30210 430
rect 30326 400 31218 430
rect 31334 400 31890 430
rect 32006 400 32898 430
rect 33014 400 33906 430
rect 34022 400 34578 430
rect 34694 400 35586 430
rect 35702 400 36594 430
rect 36710 400 37266 430
rect 37382 400 38274 430
rect 38390 400 39282 430
rect 39398 400 39954 430
rect 40070 400 40962 430
rect 41078 400 41970 430
rect 42086 400 42642 430
rect 42758 400 43650 430
rect 43766 400 44658 430
rect 44774 400 45330 430
rect 45446 400 46338 430
rect 46454 400 47346 430
rect 47462 400 48018 430
rect 48134 400 49026 430
rect 49142 400 50034 430
rect 50150 400 50706 430
rect 50822 400 51714 430
rect 51830 400 52722 430
rect 52838 400 53394 430
rect 53510 400 54402 430
rect 54518 400 55410 430
rect 55526 400 56082 430
rect 56198 400 57090 430
rect 57206 400 58098 430
rect 58214 400 58770 430
rect 58886 400 59778 430
rect 59894 400 60786 430
rect 60902 400 61458 430
rect 61574 400 62466 430
rect 62582 400 63474 430
rect 63590 400 64146 430
rect 64262 400 65154 430
rect 65270 400 66162 430
rect 66278 400 66834 430
rect 66950 400 67842 430
rect 67958 400 68850 430
rect 68966 400 69522 430
rect 69638 400 70530 430
rect 70646 400 71538 430
rect 71654 400 72210 430
rect 72326 400 73218 430
rect 73334 400 74226 430
rect 74342 400 74898 430
rect 75014 400 75906 430
rect 76022 400 76914 430
rect 77030 400 77586 430
<< metal3 >>
rect 100 107184 400 107240
rect 77600 107184 77900 107240
rect 100 106176 400 106232
rect 77600 106176 77900 106232
rect 100 105504 400 105560
rect 77600 105504 77900 105560
rect 100 104496 400 104552
rect 77600 104496 77900 104552
rect 100 103488 400 103544
rect 77600 103488 77900 103544
rect 100 102816 400 102872
rect 77600 102816 77900 102872
rect 100 101808 400 101864
rect 77600 101808 77900 101864
rect 100 100800 400 100856
rect 77600 100800 77900 100856
rect 100 100128 400 100184
rect 77600 100128 77900 100184
rect 100 99120 400 99176
rect 77600 99120 77900 99176
rect 100 98112 400 98168
rect 77600 98112 77900 98168
rect 100 97440 400 97496
rect 77600 97440 77900 97496
rect 100 96432 400 96488
rect 77600 96432 77900 96488
rect 100 95424 400 95480
rect 77600 95424 77900 95480
rect 100 94752 400 94808
rect 77600 94752 77900 94808
rect 100 93744 400 93800
rect 77600 93744 77900 93800
rect 100 92736 400 92792
rect 77600 92736 77900 92792
rect 100 92064 400 92120
rect 77600 92064 77900 92120
rect 100 91056 400 91112
rect 77600 91056 77900 91112
rect 100 90384 400 90440
rect 77600 90048 77900 90104
rect 100 89376 400 89432
rect 77600 89376 77900 89432
rect 100 88368 400 88424
rect 77600 88368 77900 88424
rect 100 87696 400 87752
rect 77600 87360 77900 87416
rect 100 86688 400 86744
rect 77600 86688 77900 86744
rect 100 85680 400 85736
rect 77600 85680 77900 85736
rect 100 85008 400 85064
rect 77600 84672 77900 84728
rect 100 84000 400 84056
rect 77600 84000 77900 84056
rect 100 82992 400 83048
rect 77600 82992 77900 83048
rect 100 82320 400 82376
rect 77600 81984 77900 82040
rect 100 81312 400 81368
rect 77600 81312 77900 81368
rect 100 80304 400 80360
rect 77600 80304 77900 80360
rect 100 79632 400 79688
rect 77600 79296 77900 79352
rect 100 78624 400 78680
rect 77600 78624 77900 78680
rect 100 77616 400 77672
rect 77600 77616 77900 77672
rect 100 76944 400 77000
rect 77600 76608 77900 76664
rect 100 75936 400 75992
rect 77600 75936 77900 75992
rect 100 74928 400 74984
rect 77600 74928 77900 74984
rect 100 74256 400 74312
rect 77600 73920 77900 73976
rect 100 73248 400 73304
rect 77600 73248 77900 73304
rect 100 72240 400 72296
rect 77600 72240 77900 72296
rect 100 71568 400 71624
rect 77600 71232 77900 71288
rect 100 70560 400 70616
rect 77600 70560 77900 70616
rect 100 69552 400 69608
rect 77600 69552 77900 69608
rect 100 68880 400 68936
rect 77600 68544 77900 68600
rect 100 67872 400 67928
rect 77600 67872 77900 67928
rect 100 66864 400 66920
rect 77600 66864 77900 66920
rect 100 66192 400 66248
rect 77600 65856 77900 65912
rect 100 65184 400 65240
rect 77600 65184 77900 65240
rect 100 64176 400 64232
rect 77600 64176 77900 64232
rect 100 63504 400 63560
rect 77600 63168 77900 63224
rect 100 62496 400 62552
rect 77600 62496 77900 62552
rect 100 61488 400 61544
rect 77600 61488 77900 61544
rect 100 60816 400 60872
rect 77600 60480 77900 60536
rect 100 59808 400 59864
rect 77600 59808 77900 59864
rect 100 58800 400 58856
rect 77600 58800 77900 58856
rect 100 58128 400 58184
rect 77600 57792 77900 57848
rect 100 57120 400 57176
rect 77600 57120 77900 57176
rect 100 56112 400 56168
rect 77600 56112 77900 56168
rect 100 55440 400 55496
rect 77600 55104 77900 55160
rect 100 54432 400 54488
rect 77600 54432 77900 54488
rect 100 53424 400 53480
rect 77600 53424 77900 53480
rect 100 52752 400 52808
rect 77600 52416 77900 52472
rect 100 51744 400 51800
rect 77600 51744 77900 51800
rect 100 50736 400 50792
rect 77600 50736 77900 50792
rect 100 50064 400 50120
rect 77600 49728 77900 49784
rect 100 49056 400 49112
rect 77600 49056 77900 49112
rect 100 48048 400 48104
rect 77600 48048 77900 48104
rect 100 47376 400 47432
rect 77600 47040 77900 47096
rect 100 46368 400 46424
rect 77600 46368 77900 46424
rect 100 45360 400 45416
rect 77600 45360 77900 45416
rect 100 44688 400 44744
rect 77600 44352 77900 44408
rect 100 43680 400 43736
rect 77600 43680 77900 43736
rect 100 42672 400 42728
rect 77600 42672 77900 42728
rect 100 42000 400 42056
rect 77600 41664 77900 41720
rect 100 40992 400 41048
rect 77600 40992 77900 41048
rect 100 39984 400 40040
rect 77600 39984 77900 40040
rect 100 39312 400 39368
rect 77600 38976 77900 39032
rect 100 38304 400 38360
rect 77600 38304 77900 38360
rect 100 37296 400 37352
rect 77600 37296 77900 37352
rect 100 36624 400 36680
rect 77600 36288 77900 36344
rect 100 35616 400 35672
rect 77600 35616 77900 35672
rect 100 34608 400 34664
rect 77600 34608 77900 34664
rect 100 33936 400 33992
rect 77600 33600 77900 33656
rect 100 32928 400 32984
rect 77600 32928 77900 32984
rect 100 31920 400 31976
rect 77600 31920 77900 31976
rect 100 31248 400 31304
rect 77600 30912 77900 30968
rect 100 30240 400 30296
rect 77600 30240 77900 30296
rect 100 29232 400 29288
rect 77600 29232 77900 29288
rect 100 28560 400 28616
rect 77600 28224 77900 28280
rect 100 27552 400 27608
rect 77600 27552 77900 27608
rect 100 26544 400 26600
rect 77600 26544 77900 26600
rect 100 25872 400 25928
rect 77600 25536 77900 25592
rect 100 24864 400 24920
rect 77600 24864 77900 24920
rect 100 23856 400 23912
rect 77600 23856 77900 23912
rect 100 23184 400 23240
rect 77600 22848 77900 22904
rect 100 22176 400 22232
rect 77600 22176 77900 22232
rect 100 21168 400 21224
rect 77600 21168 77900 21224
rect 100 20496 400 20552
rect 77600 20160 77900 20216
rect 100 19488 400 19544
rect 77600 19488 77900 19544
rect 100 18480 400 18536
rect 77600 18480 77900 18536
rect 100 17808 400 17864
rect 77600 17472 77900 17528
rect 100 16800 400 16856
rect 77600 16800 77900 16856
rect 100 15792 400 15848
rect 77600 15792 77900 15848
rect 100 15120 400 15176
rect 77600 15120 77900 15176
rect 100 14112 400 14168
rect 77600 14112 77900 14168
rect 100 13104 400 13160
rect 77600 13104 77900 13160
rect 100 12432 400 12488
rect 77600 12432 77900 12488
rect 100 11424 400 11480
rect 77600 11424 77900 11480
rect 100 10416 400 10472
rect 77600 10416 77900 10472
rect 100 9744 400 9800
rect 77600 9744 77900 9800
rect 100 8736 400 8792
rect 77600 8736 77900 8792
rect 100 7728 400 7784
rect 77600 7728 77900 7784
rect 100 7056 400 7112
rect 77600 7056 77900 7112
rect 100 6048 400 6104
rect 77600 6048 77900 6104
rect 100 5040 400 5096
rect 77600 5040 77900 5096
rect 100 4368 400 4424
rect 77600 4368 77900 4424
rect 100 3360 400 3416
rect 77600 3360 77900 3416
rect 100 2352 400 2408
rect 77600 2352 77900 2408
rect 100 1680 400 1736
rect 77600 1680 77900 1736
rect 100 672 400 728
rect 77600 672 77900 728
<< obsm3 >>
rect 9 107154 70 107226
rect 430 107154 77570 107226
rect 9 106262 77658 107154
rect 9 106146 70 106262
rect 430 106146 77570 106262
rect 9 105590 77658 106146
rect 9 105474 70 105590
rect 430 105474 77570 105590
rect 9 104582 77658 105474
rect 9 104466 70 104582
rect 430 104466 77570 104582
rect 9 103574 77658 104466
rect 9 103458 70 103574
rect 430 103458 77570 103574
rect 9 102902 77658 103458
rect 9 102786 70 102902
rect 430 102786 77570 102902
rect 9 101894 77658 102786
rect 9 101778 70 101894
rect 430 101778 77570 101894
rect 9 100886 77658 101778
rect 9 100770 70 100886
rect 430 100770 77570 100886
rect 9 100214 77658 100770
rect 9 100098 70 100214
rect 430 100098 77570 100214
rect 9 99206 77658 100098
rect 9 99090 70 99206
rect 430 99090 77570 99206
rect 9 98198 77658 99090
rect 9 98082 70 98198
rect 430 98082 77570 98198
rect 9 97526 77658 98082
rect 9 97410 70 97526
rect 430 97410 77570 97526
rect 9 96518 77658 97410
rect 9 96402 70 96518
rect 430 96402 77570 96518
rect 9 95510 77658 96402
rect 9 95394 70 95510
rect 430 95394 77570 95510
rect 9 94838 77658 95394
rect 9 94722 70 94838
rect 430 94722 77570 94838
rect 9 93830 77658 94722
rect 9 93714 70 93830
rect 430 93714 77570 93830
rect 9 92822 77658 93714
rect 9 92706 70 92822
rect 430 92706 77570 92822
rect 9 92150 77658 92706
rect 9 92034 70 92150
rect 430 92034 77570 92150
rect 9 91142 77658 92034
rect 9 91026 70 91142
rect 430 91026 77570 91142
rect 9 90470 77658 91026
rect 9 90354 70 90470
rect 430 90354 77658 90470
rect 9 90134 77658 90354
rect 9 90018 77570 90134
rect 9 89462 77658 90018
rect 9 89346 70 89462
rect 430 89346 77570 89462
rect 9 88454 77658 89346
rect 9 88338 70 88454
rect 430 88338 77570 88454
rect 9 87782 77658 88338
rect 9 87666 70 87782
rect 430 87666 77658 87782
rect 9 87446 77658 87666
rect 9 87330 77570 87446
rect 9 86774 77658 87330
rect 9 86658 70 86774
rect 430 86658 77570 86774
rect 9 85766 77658 86658
rect 9 85650 70 85766
rect 430 85650 77570 85766
rect 9 85094 77658 85650
rect 9 84978 70 85094
rect 430 84978 77658 85094
rect 9 84758 77658 84978
rect 9 84642 77570 84758
rect 9 84086 77658 84642
rect 9 83970 70 84086
rect 430 83970 77570 84086
rect 9 83078 77658 83970
rect 9 82962 70 83078
rect 430 82962 77570 83078
rect 9 82406 77658 82962
rect 9 82290 70 82406
rect 430 82290 77658 82406
rect 9 82070 77658 82290
rect 9 81954 77570 82070
rect 9 81398 77658 81954
rect 9 81282 70 81398
rect 430 81282 77570 81398
rect 9 80390 77658 81282
rect 9 80274 70 80390
rect 430 80274 77570 80390
rect 9 79718 77658 80274
rect 9 79602 70 79718
rect 430 79602 77658 79718
rect 9 79382 77658 79602
rect 9 79266 77570 79382
rect 9 78710 77658 79266
rect 9 78594 70 78710
rect 430 78594 77570 78710
rect 9 77702 77658 78594
rect 9 77586 70 77702
rect 430 77586 77570 77702
rect 9 77030 77658 77586
rect 9 76914 70 77030
rect 430 76914 77658 77030
rect 9 76694 77658 76914
rect 9 76578 77570 76694
rect 9 76022 77658 76578
rect 9 75906 70 76022
rect 430 75906 77570 76022
rect 9 75014 77658 75906
rect 9 74898 70 75014
rect 430 74898 77570 75014
rect 9 74342 77658 74898
rect 9 74226 70 74342
rect 430 74226 77658 74342
rect 9 74006 77658 74226
rect 9 73890 77570 74006
rect 9 73334 77658 73890
rect 9 73218 70 73334
rect 430 73218 77570 73334
rect 9 72326 77658 73218
rect 9 72210 70 72326
rect 430 72210 77570 72326
rect 9 71654 77658 72210
rect 9 71538 70 71654
rect 430 71538 77658 71654
rect 9 71318 77658 71538
rect 9 71202 77570 71318
rect 9 70646 77658 71202
rect 9 70530 70 70646
rect 430 70530 77570 70646
rect 9 69638 77658 70530
rect 9 69522 70 69638
rect 430 69522 77570 69638
rect 9 68966 77658 69522
rect 9 68850 70 68966
rect 430 68850 77658 68966
rect 9 68630 77658 68850
rect 9 68514 77570 68630
rect 9 67958 77658 68514
rect 9 67842 70 67958
rect 430 67842 77570 67958
rect 9 66950 77658 67842
rect 9 66834 70 66950
rect 430 66834 77570 66950
rect 9 66278 77658 66834
rect 9 66162 70 66278
rect 430 66162 77658 66278
rect 9 65942 77658 66162
rect 9 65826 77570 65942
rect 9 65270 77658 65826
rect 9 65154 70 65270
rect 430 65154 77570 65270
rect 9 64262 77658 65154
rect 9 64146 70 64262
rect 430 64146 77570 64262
rect 9 63590 77658 64146
rect 9 63474 70 63590
rect 430 63474 77658 63590
rect 9 63254 77658 63474
rect 9 63138 77570 63254
rect 9 62582 77658 63138
rect 9 62466 70 62582
rect 430 62466 77570 62582
rect 9 61574 77658 62466
rect 9 61458 70 61574
rect 430 61458 77570 61574
rect 9 60902 77658 61458
rect 9 60786 70 60902
rect 430 60786 77658 60902
rect 9 60566 77658 60786
rect 9 60450 77570 60566
rect 9 59894 77658 60450
rect 9 59778 70 59894
rect 430 59778 77570 59894
rect 9 58886 77658 59778
rect 9 58770 70 58886
rect 430 58770 77570 58886
rect 9 58214 77658 58770
rect 9 58098 70 58214
rect 430 58098 77658 58214
rect 9 57878 77658 58098
rect 9 57762 77570 57878
rect 9 57206 77658 57762
rect 9 57090 70 57206
rect 430 57090 77570 57206
rect 9 56198 77658 57090
rect 9 56082 70 56198
rect 430 56082 77570 56198
rect 9 55526 77658 56082
rect 9 55410 70 55526
rect 430 55410 77658 55526
rect 9 55190 77658 55410
rect 9 55074 77570 55190
rect 9 54518 77658 55074
rect 9 54402 70 54518
rect 430 54402 77570 54518
rect 9 53510 77658 54402
rect 9 53394 70 53510
rect 430 53394 77570 53510
rect 9 52838 77658 53394
rect 9 52722 70 52838
rect 430 52722 77658 52838
rect 9 52502 77658 52722
rect 9 52386 77570 52502
rect 9 51830 77658 52386
rect 9 51714 70 51830
rect 430 51714 77570 51830
rect 9 50822 77658 51714
rect 9 50706 70 50822
rect 430 50706 77570 50822
rect 9 50150 77658 50706
rect 9 50034 70 50150
rect 430 50034 77658 50150
rect 9 49814 77658 50034
rect 9 49698 77570 49814
rect 9 49142 77658 49698
rect 9 49026 70 49142
rect 430 49026 77570 49142
rect 9 48134 77658 49026
rect 9 48018 70 48134
rect 430 48018 77570 48134
rect 9 47462 77658 48018
rect 9 47346 70 47462
rect 430 47346 77658 47462
rect 9 47126 77658 47346
rect 9 47010 77570 47126
rect 9 46454 77658 47010
rect 9 46338 70 46454
rect 430 46338 77570 46454
rect 9 45446 77658 46338
rect 9 45330 70 45446
rect 430 45330 77570 45446
rect 9 44774 77658 45330
rect 9 44658 70 44774
rect 430 44658 77658 44774
rect 9 44438 77658 44658
rect 9 44322 77570 44438
rect 9 43766 77658 44322
rect 9 43650 70 43766
rect 430 43650 77570 43766
rect 9 42758 77658 43650
rect 9 42642 70 42758
rect 430 42642 77570 42758
rect 9 42086 77658 42642
rect 9 41970 70 42086
rect 430 41970 77658 42086
rect 9 41750 77658 41970
rect 9 41634 77570 41750
rect 9 41078 77658 41634
rect 9 40962 70 41078
rect 430 40962 77570 41078
rect 9 40070 77658 40962
rect 9 39954 70 40070
rect 430 39954 77570 40070
rect 9 39398 77658 39954
rect 9 39282 70 39398
rect 430 39282 77658 39398
rect 9 39062 77658 39282
rect 9 38946 77570 39062
rect 9 38390 77658 38946
rect 9 38274 70 38390
rect 430 38274 77570 38390
rect 9 37382 77658 38274
rect 9 37266 70 37382
rect 430 37266 77570 37382
rect 9 36710 77658 37266
rect 9 36594 70 36710
rect 430 36594 77658 36710
rect 9 36374 77658 36594
rect 9 36258 77570 36374
rect 9 35702 77658 36258
rect 9 35586 70 35702
rect 430 35586 77570 35702
rect 9 34694 77658 35586
rect 9 34578 70 34694
rect 430 34578 77570 34694
rect 9 34022 77658 34578
rect 9 33906 70 34022
rect 430 33906 77658 34022
rect 9 33686 77658 33906
rect 9 33570 77570 33686
rect 9 33014 77658 33570
rect 9 32898 70 33014
rect 430 32898 77570 33014
rect 9 32006 77658 32898
rect 9 31890 70 32006
rect 430 31890 77570 32006
rect 9 31334 77658 31890
rect 9 31218 70 31334
rect 430 31218 77658 31334
rect 9 30998 77658 31218
rect 9 30882 77570 30998
rect 9 30326 77658 30882
rect 9 30210 70 30326
rect 430 30210 77570 30326
rect 9 29318 77658 30210
rect 9 29202 70 29318
rect 430 29202 77570 29318
rect 9 28646 77658 29202
rect 9 28530 70 28646
rect 430 28530 77658 28646
rect 9 28310 77658 28530
rect 9 28194 77570 28310
rect 9 27638 77658 28194
rect 9 27522 70 27638
rect 430 27522 77570 27638
rect 9 26630 77658 27522
rect 9 26514 70 26630
rect 430 26514 77570 26630
rect 9 25958 77658 26514
rect 9 25842 70 25958
rect 430 25842 77658 25958
rect 9 25622 77658 25842
rect 9 25506 77570 25622
rect 9 24950 77658 25506
rect 9 24834 70 24950
rect 430 24834 77570 24950
rect 9 23942 77658 24834
rect 9 23826 70 23942
rect 430 23826 77570 23942
rect 9 23270 77658 23826
rect 9 23154 70 23270
rect 430 23154 77658 23270
rect 9 22934 77658 23154
rect 9 22818 77570 22934
rect 9 22262 77658 22818
rect 9 22146 70 22262
rect 430 22146 77570 22262
rect 9 21254 77658 22146
rect 9 21138 70 21254
rect 430 21138 77570 21254
rect 9 20582 77658 21138
rect 9 20466 70 20582
rect 430 20466 77658 20582
rect 9 20246 77658 20466
rect 9 20130 77570 20246
rect 9 19574 77658 20130
rect 9 19458 70 19574
rect 430 19458 77570 19574
rect 9 18566 77658 19458
rect 9 18450 70 18566
rect 430 18450 77570 18566
rect 9 17894 77658 18450
rect 9 17778 70 17894
rect 430 17778 77658 17894
rect 9 17558 77658 17778
rect 9 17442 77570 17558
rect 9 16886 77658 17442
rect 9 16770 70 16886
rect 430 16770 77570 16886
rect 9 15878 77658 16770
rect 9 15762 70 15878
rect 430 15762 77570 15878
rect 9 15206 77658 15762
rect 9 15090 70 15206
rect 430 15090 77570 15206
rect 9 14198 77658 15090
rect 9 14082 70 14198
rect 430 14082 77570 14198
rect 9 13190 77658 14082
rect 9 13074 70 13190
rect 430 13074 77570 13190
rect 9 12518 77658 13074
rect 9 12402 70 12518
rect 430 12402 77570 12518
rect 9 11510 77658 12402
rect 9 11394 70 11510
rect 430 11394 77570 11510
rect 9 10502 77658 11394
rect 9 10386 70 10502
rect 430 10386 77570 10502
rect 9 9830 77658 10386
rect 9 9714 70 9830
rect 430 9714 77570 9830
rect 9 8822 77658 9714
rect 9 8706 70 8822
rect 430 8706 77570 8822
rect 9 7814 77658 8706
rect 9 7698 70 7814
rect 430 7698 77570 7814
rect 9 7142 77658 7698
rect 9 7026 70 7142
rect 430 7026 77570 7142
rect 9 6134 77658 7026
rect 9 6018 70 6134
rect 430 6018 77570 6134
rect 9 5126 77658 6018
rect 9 5010 70 5126
rect 430 5010 77570 5126
rect 9 4454 77658 5010
rect 9 4338 70 4454
rect 430 4338 77570 4454
rect 9 3446 77658 4338
rect 9 3330 70 3446
rect 430 3330 77570 3446
rect 9 2438 77658 3330
rect 9 2322 70 2438
rect 430 2322 77570 2438
rect 9 1766 77658 2322
rect 9 1650 70 1766
rect 430 1650 77570 1766
rect 9 798 77658 1650
<< metal4 >>
rect 2224 1538 2384 106262
rect 9904 1538 10064 106262
rect 17584 1538 17744 106262
rect 25264 1538 25424 106262
rect 32944 1538 33104 106262
rect 40624 1538 40784 106262
rect 48304 1538 48464 106262
rect 55984 1538 56144 106262
rect 63664 1538 63824 106262
rect 71344 1538 71504 106262
<< obsm4 >>
rect 1666 11601 2194 92447
rect 2414 11601 9874 92447
rect 10094 11601 17554 92447
rect 17774 11601 25234 92447
rect 25454 11601 32914 92447
rect 33134 11601 40594 92447
rect 40814 11601 48274 92447
rect 48494 11601 55954 92447
rect 56174 11601 63634 92447
rect 63854 11601 68810 92447
<< labels >>
rlabel metal3 s 100 64176 400 64232 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 65184 400 65240 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 31920 400 31976 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 56112 400 56168 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 38304 400 38360 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 32928 400 32984 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 33936 107600 33992 107900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 77600 33600 77900 33656 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 77600 102816 77900 102872 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47376 107600 47432 107900 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 77600 13104 77900 13160 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 100 104496 400 104552 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 59136 107600 59192 107900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 65184 100 65240 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 77616 107600 77672 107900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 77600 95424 77900 95480 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 76944 100 77000 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 12432 100 12488 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 77616 400 77672 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 63504 400 63560 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 72240 400 72296 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 58128 400 58184 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 77600 107184 77900 107240 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 60816 100 60872 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 77600 672 77900 728 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 9744 400 9800 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 100 82992 400 83048 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 67872 107600 67928 107900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 77600 97440 77900 97496 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 77600 85680 77900 85736 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 77600 106176 77900 106232 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 77600 57120 77900 57176 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 17808 400 17864 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 77600 32928 77900 32984 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 60816 107600 60872 107900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 42672 400 42728 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 48048 400 48104 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 77600 80304 77900 80360 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 77600 74928 77900 74984 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 100 96432 400 96488 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 57120 100 57176 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 23856 400 23912 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 77600 7056 77900 7112 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 43680 107600 43736 107900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 26544 100 26600 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 8736 100 8792 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 97440 400 97496 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 17808 107600 17864 107900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9744 107600 9800 107900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 38304 107600 38360 107900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 77600 1680 77900 1736 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 77600 38976 77900 39032 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 75264 107600 75320 107900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 26544 400 26600 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 13104 400 13160 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 100 85008 400 85064 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 77616 100 77672 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 100 94752 400 94808 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 77600 62496 77900 62552 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 77600 50736 77900 50792 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 77600 9744 77900 9800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 28560 400 28616 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 66192 107600 66248 107900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 77600 30240 77900 30296 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 75936 400 75992 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 77600 99120 77900 99176 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 36624 107600 36680 107900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 77600 52416 77900 52472 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 69552 400 69608 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 12432 400 12488 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 52752 107600 52808 107900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 73248 400 73304 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 29568 107600 29624 107900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 46368 400 46424 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 77600 105504 77900 105560 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 0 107600 56 107900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 13440 107600 13496 107900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 59808 100 59864 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 75936 107600 75992 107900 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 92736 400 92792 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 68880 400 68936 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37296 100 37352 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 77600 92736 77900 92792 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 10416 100 10472 400 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 77600 8736 77900 8792 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 5376 107600 5432 107900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6048 100 6104 400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 77600 23856 77900 23912 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 61488 400 61544 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 77600 35616 77900 35672 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 34608 400 34664 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 77600 3360 77900 3416 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 77600 17472 77900 17528 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 39312 100 39368 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 31248 100 31304 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 50064 107600 50120 107900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 63504 100 63560 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 77600 48048 77900 48104 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 69888 107600 69944 107900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 32928 100 32984 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 43008 107600 43064 107900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 33936 400 33992 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 61488 100 61544 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 55440 100 55496 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 22176 100 22232 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 4368 400 4424 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 27552 107600 27608 107900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 42672 100 42728 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24192 107600 24248 107900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 16800 400 16856 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 52752 400 52808 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 67872 100 67928 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23856 100 23912 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 77600 101808 77900 101864 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 77600 56112 77900 56168 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 28560 100 28616 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 22176 107600 22232 107900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 100 81312 400 81368 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 77600 81984 77900 82040 6 la_data_in[15]
port 121 nsew signal input
rlabel metal3 s 100 101808 400 101864 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 77600 29232 77900 29288 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 31248 107600 31304 107900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 14112 400 14168 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 6048 107600 6104 107900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 77600 34608 77900 34664 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 70560 400 70616 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 40992 400 41048 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 77600 84672 77900 84728 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 32256 107600 32312 107900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 4368 107600 4424 107900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 42000 107600 42056 107900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 100 84000 400 84056 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 87696 400 87752 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 77600 38304 77900 38360 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 25872 107600 25928 107900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 7056 400 7112 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 63504 107600 63560 107900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 37296 400 37352 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 62496 400 62552 6 la_data_in[33]
port 141 nsew signal input
rlabel metal3 s 100 100128 400 100184 6 la_data_in[34]
port 142 nsew signal input
rlabel metal3 s 100 82320 400 82376 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 66192 100 66248 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal3 s 100 91056 400 91112 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 42000 100 42056 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 35616 107600 35672 107900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 77600 65856 77900 65912 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 31920 100 31976 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 44688 100 44744 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 31248 400 31304 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 72576 107600 72632 107900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 77600 15792 77900 15848 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 30240 100 30296 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 77600 82992 77900 83048 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 58128 100 58184 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 28560 107600 28616 107900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 20496 107600 20552 107900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal3 s 100 100800 400 100856 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 21504 107600 21560 107900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 43680 100 43736 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 77600 46368 77900 46424 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 57120 107600 57176 107900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 51072 107600 51128 107900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 27552 400 27608 6 la_data_in[56]
port 166 nsew signal input
rlabel metal3 s 100 95424 400 95480 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 33936 100 33992 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 77600 100128 77900 100184 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 15792 100 15848 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 77600 76608 77900 76664 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 2352 400 2408 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 54432 100 54488 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 8736 107600 8792 107900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 18480 100 18536 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 77600 49056 77900 49112 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1680 400 1736 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 68880 107600 68936 107900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 65184 107600 65240 107900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 77600 65184 77900 65240 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 3360 400 3416 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 66864 400 66920 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 34608 100 34664 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 77600 53424 77900 53480 6 la_data_out[14]
port 184 nsew signal output
rlabel metal3 s 100 79632 400 79688 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 77600 66864 77900 66920 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 30240 107600 30296 107900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 77600 92064 77900 92120 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 49056 100 49112 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 77600 58800 77900 58856 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 77600 28224 77900 28280 6 la_data_out[20]
port 191 nsew signal output
rlabel metal3 s 100 92064 400 92120 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 77600 73248 77900 73304 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 27552 100 27608 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 42000 400 42056 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 50064 100 50120 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 90384 400 90440 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 40992 107600 41048 107900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 77600 89376 77900 89432 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 39984 100 40040 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 21168 400 21224 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 77600 57792 77900 57848 6 la_data_out[30]
port 202 nsew signal output
rlabel metal3 s 77600 19488 77900 19544 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 39312 107600 39368 107900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 77600 31920 77900 31976 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 45360 100 45416 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 34944 107600 35000 107900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 77600 90048 77900 90104 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 77600 51744 77900 51800 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 77600 16800 77900 16856 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 77600 27552 77900 27608 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 15120 400 15176 6 la_data_out[3]
port 212 nsew signal output
rlabel metal3 s 77600 12432 77900 12488 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 77600 43680 77900 43736 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 77600 93744 77900 93800 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 5040 100 5096 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 38304 100 38360 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal3 s 100 107184 400 107240 6 la_data_out[45]
port 218 nsew signal output
rlabel metal3 s 100 106176 400 106232 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 66192 400 66248 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 21168 100 21224 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal3 s 77600 6048 77900 6104 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 37632 107600 37688 107900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 16800 107600 16856 107900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal3 s 100 89376 400 89432 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 77600 21168 77900 21224 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 88368 400 88424 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 77600 78624 77900 78680 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 19488 107600 19544 107900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 77600 37296 77900 37352 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 55440 107600 55496 107900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 77600 79296 77900 79352 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 35616 400 35672 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 77600 70560 77900 70616 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 59808 107600 59864 107900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 24864 100 24920 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal3 s 77600 2352 77900 2408 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 77600 22176 77900 22232 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 77600 41664 77900 41720 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 74256 107600 74312 107900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 5040 400 5096 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 77600 59808 77900 59864 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 77600 49728 77900 49784 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 77600 81312 77900 81368 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 77600 67872 77900 67928 6 la_oenb[11]
port 245 nsew signal input
rlabel metal3 s 100 93744 400 93800 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 74256 400 74312 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 68880 100 68936 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal3 s 77600 4368 77900 4424 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 13104 100 13160 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 11424 400 11480 6 la_oenb[17]
port 251 nsew signal input
rlabel metal3 s 100 99120 400 99176 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 77600 22848 77900 22904 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 2688 107600 2744 107900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 23184 107600 23240 107900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 53760 107600 53816 107900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 25872 100 25928 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 77600 72240 77900 72296 6 la_oenb[24]
port 259 nsew signal input
rlabel metal3 s 77600 5040 77900 5096 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 3360 107600 3416 107900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 16800 100 16856 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 57120 400 57176 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 77600 103488 77900 103544 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 76944 107600 77000 107900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 77600 94752 77900 94808 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 24864 107600 24920 107900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 77600 91056 77900 91112 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 47376 100 47432 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 672 107600 728 107900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 2352 100 2408 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 672 100 728 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal3 s 100 105504 400 105560 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 48048 100 48104 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 39984 400 40040 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 50736 400 50792 6 la_oenb[3]
port 276 nsew signal input
rlabel metal3 s 77600 26544 77900 26600 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 18816 107600 18872 107900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 58800 400 58856 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 17808 100 17864 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 40992 100 41048 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 61824 107600 61880 107900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 74256 100 74312 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 10416 400 10472 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 67872 400 67928 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 672 400 728 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 100 86688 400 86744 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 71568 100 71624 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 15120 107600 15176 107900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal3 s 77600 14112 77900 14168 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 77600 73920 77900 73976 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 50064 400 50120 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 77600 63168 77900 63224 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 70560 100 70616 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 67200 107600 67256 107900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal3 s 77600 24864 77900 24920 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 40320 107600 40376 107900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal3 s 77600 7728 77900 7784 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 45360 400 45416 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 11424 100 11480 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 77600 61488 77900 61544 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 22176 400 22232 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 77600 75936 77900 75992 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 23184 100 23240 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal3 s 77600 10416 77900 10472 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 11424 107600 11480 107900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 64512 107600 64568 107900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 77600 86688 77900 86744 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 8064 107600 8120 107900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 59808 400 59864 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 106262 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 106262 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 106262 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 106262 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 106262 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 106262 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 106262 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 106262 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 106262 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 106262 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 77600 30912 77900 30968 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 1680 107600 1736 107900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 77600 47040 77900 47096 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 46368 107600 46424 107900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 26880 107600 26936 107900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 53424 400 53480 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 7728 100 7784 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 51744 100 51800 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 8736 400 8792 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 77600 77616 77900 77672 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 58800 100 58856 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 51744 400 51800 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 77600 44352 77900 44408 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 77600 11424 77900 11480 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 6048 400 6104 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 71568 107600 71624 107900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 52752 100 52808 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 74928 100 74984 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 77600 36288 77900 36344 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal3 s 100 103488 400 103544 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 15792 400 15848 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 16128 107600 16184 107900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 77600 69552 77900 69608 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 77600 104496 77900 104552 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 36624 100 36680 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 36624 400 36680 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 77600 54432 77900 54488 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 72240 100 72296 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 56448 107600 56504 107900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 69552 100 69608 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 23184 400 23240 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 4368 100 4424 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal3 s 77600 15120 77900 15176 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 77600 39984 77900 40040 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 14112 107600 14168 107900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 77600 96432 77900 96488 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 71568 400 71624 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal3 s 100 78624 400 78680 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 74928 400 74984 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 3360 100 3416 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 19488 400 19544 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 77600 64176 77900 64232 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 53424 100 53480 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 48384 107600 48440 107900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 70560 107600 70616 107900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal3 s 100 98112 400 98168 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 14112 100 14168 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 73248 107600 73304 107900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 55440 400 55496 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 77600 88368 77900 88424 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 77600 45360 77900 45416 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 64176 100 64232 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 62496 107600 62552 107900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 7056 107600 7112 107900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 29232 100 29288 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 77600 71232 77900 71288 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 75936 100 75992 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 77600 42672 77900 42728 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 49056 400 49112 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal3 s 77600 18480 77900 18536 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 15120 100 15176 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 46368 100 46424 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 77600 55104 77900 55160 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 58128 107600 58184 107900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 77600 98112 77900 98168 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal3 s 77600 20160 77900 20216 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 18480 400 18536 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 77600 68544 77900 68600 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1680 100 1736 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 77600 100800 77900 100856 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 54432 107600 54488 107900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal3 s 77600 25536 77900 25592 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 51744 107600 51800 107900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 25872 400 25928 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 29232 400 29288 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 62496 100 62552 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 73248 100 73304 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 44688 400 44744 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal3 s 100 80304 400 80360 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 10752 107600 10808 107900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 30240 400 30296 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 19488 100 19544 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 7056 100 7112 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 32928 107600 32984 107900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 12432 107600 12488 107900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 50736 100 50792 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 49056 107600 49112 107900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 77600 40992 77900 41048 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 60816 400 60872 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 77600 87360 77900 87416 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 20496 100 20552 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 35616 100 35672 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 7728 400 7784 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 77600 84000 77900 84056 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 56112 100 56168 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 45696 107600 45752 107900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 44688 107600 44744 107900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal3 s 100 85680 400 85736 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal3 s 100 102816 400 102872 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 66864 100 66920 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 20496 400 20552 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 76944 400 77000 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 77600 60480 77900 60536 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 78000 108000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 19749118
string GDS_FILE /home/runner/work/gf0mpw-serv-array/gf0mpw-serv-array/openlane/tiny_user_project/runs/22_12_02_14_26/results/signoff/tiny_user_project.magic.gds
string GDS_START 294472
<< end >>

