magic
tech gf180mcuC
magscale 1 5
timestamp 1670250507
<< obsm1 >>
rect 672 1538 99288 58438
<< obsm2 >>
rect 2238 1465 99218 58427
<< metal3 >>
rect 99800 57792 100000 57848
rect 99800 53816 100000 53872
rect 99800 49840 100000 49896
rect 99800 45864 100000 45920
rect 99800 41888 100000 41944
rect 99800 37912 100000 37968
rect 99800 33936 100000 33992
rect 99800 29960 100000 30016
rect 99800 25984 100000 26040
rect 99800 22008 100000 22064
rect 99800 18032 100000 18088
rect 99800 14056 100000 14112
rect 99800 10080 100000 10136
rect 99800 6104 100000 6160
rect 99800 2128 100000 2184
<< obsm3 >>
rect 2233 57878 99800 58422
rect 2233 57762 99770 57878
rect 2233 53902 99800 57762
rect 2233 53786 99770 53902
rect 2233 49926 99800 53786
rect 2233 49810 99770 49926
rect 2233 45950 99800 49810
rect 2233 45834 99770 45950
rect 2233 41974 99800 45834
rect 2233 41858 99770 41974
rect 2233 37998 99800 41858
rect 2233 37882 99770 37998
rect 2233 34022 99800 37882
rect 2233 33906 99770 34022
rect 2233 30046 99800 33906
rect 2233 29930 99770 30046
rect 2233 26070 99800 29930
rect 2233 25954 99770 26070
rect 2233 22094 99800 25954
rect 2233 21978 99770 22094
rect 2233 18118 99800 21978
rect 2233 18002 99770 18118
rect 2233 14142 99800 18002
rect 2233 14026 99770 14142
rect 2233 10166 99800 14026
rect 2233 10050 99770 10166
rect 2233 6190 99800 10050
rect 2233 6074 99770 6190
rect 2233 2214 99800 6074
rect 2233 2098 99770 2214
rect 2233 1470 99800 2098
<< metal4 >>
rect 2224 1538 2384 58438
rect 4474 1538 4634 58438
rect 6724 1538 6884 58438
rect 8974 1538 9134 58438
rect 11224 1538 11384 58438
rect 13474 1538 13634 58438
rect 15724 1538 15884 58438
rect 17974 1538 18134 58438
rect 20224 1538 20384 58438
rect 22474 1538 22634 58438
rect 24724 1538 24884 58438
rect 26974 1538 27134 58438
rect 29224 1538 29384 58438
rect 31474 1538 31634 58438
rect 33724 1538 33884 58438
rect 35974 1538 36134 58438
rect 38224 1538 38384 58438
rect 40474 1538 40634 58438
rect 42724 1538 42884 58438
rect 44974 1538 45134 58438
rect 47224 1538 47384 58438
rect 49474 1538 49634 58438
rect 51724 1538 51884 58438
rect 53974 1538 54134 58438
rect 56224 1538 56384 58438
rect 58474 1538 58634 58438
rect 60724 1538 60884 58438
rect 62974 1538 63134 58438
rect 65224 1538 65384 58438
rect 67474 1538 67634 58438
rect 69724 1538 69884 58438
rect 71974 1538 72134 58438
rect 74224 1538 74384 58438
rect 76474 1538 76634 58438
rect 78724 1538 78884 58438
rect 80974 1538 81134 58438
rect 83224 1538 83384 58438
rect 85474 1538 85634 58438
rect 87724 1538 87884 58438
rect 89974 1538 90134 58438
rect 92224 1538 92384 58438
rect 94474 1538 94634 58438
rect 96724 1538 96884 58438
rect 98974 1538 99134 58438
<< obsm4 >>
rect 39438 1508 40444 27767
rect 40664 1508 42694 27767
rect 42914 1508 44944 27767
rect 45164 1508 47194 27767
rect 47414 1508 49444 27767
rect 49664 1508 51694 27767
rect 51914 1508 53944 27767
rect 54164 1508 56194 27767
rect 56414 1508 58444 27767
rect 58664 1508 60694 27767
rect 60914 1508 62944 27767
rect 63164 1508 65194 27767
rect 65414 1508 67444 27767
rect 67664 1508 69694 27767
rect 69914 1508 71944 27767
rect 72164 1508 74194 27767
rect 74414 1508 76444 27767
rect 76664 1508 78694 27767
rect 78914 1508 80944 27767
rect 81164 1508 83194 27767
rect 83414 1508 85444 27767
rect 85664 1508 87694 27767
rect 87914 1508 89944 27767
rect 90164 1508 91378 27767
rect 39438 1465 91378 1508
<< labels >>
rlabel metal3 s 99800 2128 100000 2184 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 99800 6104 100000 6160 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 99800 10080 100000 10136 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 99800 14056 100000 14112 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 99800 18032 100000 18088 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 99800 41888 100000 41944 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 99800 45864 100000 45920 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 99800 49840 100000 49896 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 99800 53816 100000 53872 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 99800 57792 100000 57848 6 io_oeb[4]
port 10 nsew signal output
rlabel metal3 s 99800 22008 100000 22064 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 99800 25984 100000 26040 6 io_out[1]
port 12 nsew signal output
rlabel metal3 s 99800 29960 100000 30016 6 io_out[2]
port 13 nsew signal output
rlabel metal3 s 99800 33936 100000 33992 6 io_out[3]
port 14 nsew signal output
rlabel metal3 s 99800 37912 100000 37968 6 io_out[4]
port 15 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 6724 1538 6884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 11224 1538 11384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 15724 1538 15884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 20224 1538 20384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 24724 1538 24884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 29224 1538 29384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 33724 1538 33884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 38224 1538 38384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 42724 1538 42884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 47224 1538 47384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 51724 1538 51884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 56224 1538 56384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 60724 1538 60884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 65224 1538 65384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 69724 1538 69884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 74224 1538 74384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 78724 1538 78884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 83224 1538 83384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 87724 1538 87884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 92224 1538 92384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 96724 1538 96884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 4474 1538 4634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 8974 1538 9134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 13474 1538 13634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 17974 1538 18134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 22474 1538 22634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 26974 1538 27134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 31474 1538 31634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 35974 1538 36134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 40474 1538 40634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 44974 1538 45134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 49474 1538 49634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 53974 1538 54134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 58474 1538 58634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 62974 1538 63134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 67474 1538 67634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 71974 1538 72134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 76474 1538 76634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 80974 1538 81134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 85474 1538 85634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 89974 1538 90134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 94474 1538 94634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 98974 1538 99134 58438 6 vss
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29005104
string GDS_FILE /home/runner/work/gf180-mpw0-serv/gf180-mpw0-serv/openlane/serv_0/runs/22_12_05_14_25/results/signoff/serv_0.magic.gds
string GDS_START 22246308
<< end >>

