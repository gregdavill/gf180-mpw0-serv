// This is the unpowered netlist.
module serv_0 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_arbiter.o_wb_cpu_adr[0] ;
 wire \u_arbiter.o_wb_cpu_adr[10] ;
 wire \u_arbiter.o_wb_cpu_adr[11] ;
 wire \u_arbiter.o_wb_cpu_adr[12] ;
 wire \u_arbiter.o_wb_cpu_adr[13] ;
 wire \u_arbiter.o_wb_cpu_adr[14] ;
 wire \u_arbiter.o_wb_cpu_adr[15] ;
 wire \u_arbiter.o_wb_cpu_adr[16] ;
 wire \u_arbiter.o_wb_cpu_adr[17] ;
 wire \u_arbiter.o_wb_cpu_adr[18] ;
 wire \u_arbiter.o_wb_cpu_adr[19] ;
 wire \u_arbiter.o_wb_cpu_adr[1] ;
 wire \u_arbiter.o_wb_cpu_adr[20] ;
 wire \u_arbiter.o_wb_cpu_adr[21] ;
 wire \u_arbiter.o_wb_cpu_adr[22] ;
 wire \u_arbiter.o_wb_cpu_adr[23] ;
 wire \u_arbiter.o_wb_cpu_adr[24] ;
 wire \u_arbiter.o_wb_cpu_adr[25] ;
 wire \u_arbiter.o_wb_cpu_adr[26] ;
 wire \u_arbiter.o_wb_cpu_adr[27] ;
 wire \u_arbiter.o_wb_cpu_adr[28] ;
 wire \u_arbiter.o_wb_cpu_adr[29] ;
 wire \u_arbiter.o_wb_cpu_adr[2] ;
 wire \u_arbiter.o_wb_cpu_adr[30] ;
 wire \u_arbiter.o_wb_cpu_adr[31] ;
 wire \u_arbiter.o_wb_cpu_adr[3] ;
 wire \u_arbiter.o_wb_cpu_adr[4] ;
 wire \u_arbiter.o_wb_cpu_adr[5] ;
 wire \u_arbiter.o_wb_cpu_adr[6] ;
 wire \u_arbiter.o_wb_cpu_adr[7] ;
 wire \u_arbiter.o_wb_cpu_adr[8] ;
 wire \u_arbiter.o_wb_cpu_adr[9] ;
 wire \u_arbiter.o_wb_cpu_cyc ;
 wire \u_arbiter.o_wb_cpu_we ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.addr[0] ;
 wire \u_cpu.rf_ram.addr[1] ;
 wire \u_cpu.rf_ram.addr[2] ;
 wire \u_cpu.rf_ram.addr[3] ;
 wire \u_cpu.rf_ram.addr[4] ;
 wire \u_cpu.rf_ram.addr[5] ;
 wire \u_cpu.rf_ram.addr[6] ;
 wire \u_cpu.rf_ram.addr[7] ;
 wire \u_cpu.rf_ram.i_waddr[0] ;
 wire \u_cpu.rf_ram.i_waddr[1] ;
 wire \u_cpu.rf_ram.i_waddr[2] ;
 wire \u_cpu.rf_ram.i_waddr[3] ;
 wire \u_cpu.rf_ram.i_waddr[4] ;
 wire \u_cpu.rf_ram.i_waddr[5] ;
 wire \u_cpu.rf_ram.i_waddr[6] ;
 wire \u_cpu.rf_ram.i_waddr[7] ;
 wire \u_cpu.rf_ram.i_wdata[0] ;
 wire \u_cpu.rf_ram.i_wdata[1] ;
 wire \u_cpu.rf_ram.i_wdata[2] ;
 wire \u_cpu.rf_ram.i_wdata[3] ;
 wire \u_cpu.rf_ram.i_wdata[4] ;
 wire \u_cpu.rf_ram.i_wdata[5] ;
 wire \u_cpu.rf_ram.i_wdata[6] ;
 wire \u_cpu.rf_ram.i_wdata[7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.o_wen_req ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.clk ;
 wire \u_scanchain_local.clk_out ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.data_out_i ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1554_ (.I(\u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1555_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1556_ (.A1(\u_cpu.rf_ram_if.rcnt[2] ),
    .A2(_1036_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1557_ (.I(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1558_ (.I(_1038_),
    .Z(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1559_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1560_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1561_ (.A1(_1039_),
    .A2(_1040_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1562_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1563_ (.I(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1564_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1565_ (.A1(_1042_),
    .A2(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1566_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1567_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1568_ (.I(\u_cpu.cpu.bne_or_bge ),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1569_ (.A1(_1046_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1570_ (.A1(_1045_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1571_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_1044_),
    .A3(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1572_ (.I(\u_cpu.cpu.decode.op26 ),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1573_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1574_ (.A1(_1041_),
    .A2(\u_cpu.cpu.decode.opcode[2] ),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1575_ (.A1(_1053_),
    .A2(_1049_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1576_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(_1052_),
    .B(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1577_ (.I(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1578_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1579_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1580_ (.I(_1045_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1581_ (.A1(\u_cpu.cpu.decode.co_mem_word ),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1582_ (.A1(_1059_),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1583_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_1053_),
    .A3(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1584_ (.A1(_1058_),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1585_ (.A1(_1057_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1586_ (.A1(_1056_),
    .A2(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1587_ (.A1(_1050_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1588_ (.I(_1037_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1589_ (.I(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1590_ (.A1(_1067_),
    .A2(_1066_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1591_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_1068_),
    .B1(_1069_),
    .B2(\u_cpu.cpu.immdec.imm24_20[3] ),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1592_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_1068_),
    .B1(_1069_),
    .B2(\u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(_1070_),
    .A2(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1594_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_1065_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1595_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_1054_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1596_ (.A1(_1038_),
    .A2(_1050_),
    .A3(_1073_),
    .A4(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1597_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_1038_),
    .B(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1598_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1599_ (.A1(_1058_),
    .A2(_1077_),
    .A3(_1062_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1600_ (.A1(_1052_),
    .A2(_1078_),
    .B(_1065_),
    .C(_1067_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1601_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_1067_),
    .B1(_1069_),
    .B2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .C(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1602_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_1068_),
    .B1(_1069_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1603_ (.A1(_1076_),
    .A2(_1080_),
    .A3(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1604_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_1066_),
    .B(_1072_),
    .C(_1082_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1605_ (.I(_1068_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1606_ (.I(_1083_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1607_ (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1608_ (.I(net2),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1609_ (.A1(_1085_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1610_ (.I(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1611_ (.A1(_1084_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1612_ (.I(_1088_),
    .Z(\u_arbiter.o_wb_cpu_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1613_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_1086_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1614_ (.I(_1089_),
    .Z(\u_arbiter.o_wb_cpu_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1615_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1616_ (.I(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1617_ (.I(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1618_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1619_ (.I(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1620_ (.I(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1621_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1622_ (.A1(_1095_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1623_ (.I(_1094_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1624_ (.A1(_1098_),
    .A2(_1096_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1625_ (.A1(_1087_),
    .A2(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1626_ (.A1(_1085_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1627_ (.I(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1628_ (.I(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1629_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1630_ (.A1(_1097_),
    .A2(_1100_),
    .B(_1104_),
    .ZN(\u_arbiter.o_wb_cpu_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1631_ (.I(_1102_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1632_ (.I(_1105_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1633_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_1099_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1634_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .A2(_1103_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1635_ (.A1(_1106_),
    .A2(_1107_),
    .B(_1108_),
    .ZN(\u_arbiter.o_wb_cpu_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1636_ (.A1(_1098_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(_1096_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1637_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1638_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .A2(_1103_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1639_ (.A1(_1106_),
    .A2(_1110_),
    .B(_1111_),
    .ZN(\u_arbiter.o_wb_cpu_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1640_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _1641_ (.A1(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1642_ (.A1(_1112_),
    .A2(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1643_ (.I(_1102_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1644_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .A2(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1645_ (.A1(_1106_),
    .A2(_1114_),
    .B(_1116_),
    .ZN(\u_arbiter.o_wb_cpu_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1646_ (.A1(_1112_),
    .A2(_1113_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1647_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_1112_),
    .A3(_1113_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1648_ (.A1(_1087_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1649_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .A2(_1115_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1650_ (.A1(_1117_),
    .A2(_1119_),
    .B(_1120_),
    .ZN(\u_arbiter.o_wb_cpu_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1651_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_1118_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1652_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .A2(_1115_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1653_ (.A1(_1106_),
    .A2(_1121_),
    .B(_1122_),
    .ZN(\u_arbiter.o_wb_cpu_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1654_ (.I(_1101_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1655_ (.I(_1123_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1656_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1657_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_1113_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1658_ (.A1(_1125_),
    .A2(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1659_ (.A1(_1125_),
    .A2(_1126_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1660_ (.A1(_1127_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1661_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .A2(_1115_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1662_ (.A1(_1124_),
    .A2(_1129_),
    .B(_1130_),
    .ZN(\u_arbiter.o_wb_cpu_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1663_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_1128_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1664_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .A2(_1115_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1665_ (.A1(_1124_),
    .A2(_1131_),
    .B(_1132_),
    .ZN(\u_arbiter.o_wb_cpu_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1666_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .A2(_1103_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1667_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1668_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1669_ (.A1(_1135_),
    .A2(_1128_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1670_ (.A1(_1134_),
    .A2(_1136_),
    .B(_1105_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1671_ (.A1(_1134_),
    .A2(_1136_),
    .B(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1672_ (.A1(_1133_),
    .A2(_1138_),
    .ZN(\u_arbiter.o_wb_cpu_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1673_ (.I(_1105_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1674_ (.A1(_1134_),
    .A2(_1136_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1675_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1676_ (.A1(_1135_),
    .A2(_1125_),
    .A3(_1126_),
    .A4(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1677_ (.I(_1101_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1678_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .A2(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1679_ (.A1(_1139_),
    .A2(_1140_),
    .A3(_1142_),
    .B(_1144_),
    .ZN(\u_arbiter.o_wb_cpu_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1680_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1681_ (.A1(_1145_),
    .A2(_1142_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1682_ (.I(_1102_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1683_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1684_ (.A1(_1124_),
    .A2(_1146_),
    .B(_1148_),
    .ZN(\u_arbiter.o_wb_cpu_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1685_ (.A1(_1145_),
    .A2(_1142_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1686_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_1145_),
    .A3(_1142_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1687_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_1143_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1688_ (.A1(_1139_),
    .A2(_1149_),
    .A3(_1150_),
    .B(_1151_),
    .ZN(\u_arbiter.o_wb_cpu_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1689_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_1150_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1690_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(_1152_),
    .S(_1087_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1691_ (.I(_1153_),
    .Z(\u_arbiter.o_wb_cpu_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1692_ (.I(_1105_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1693_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_1150_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1694_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1695_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_1142_),
    .A4(_1156_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1696_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .A2(_1143_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1697_ (.A1(_1154_),
    .A2(_1155_),
    .A3(_1157_),
    .B(_1158_),
    .ZN(\u_arbiter.o_wb_cpu_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1698_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_1157_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1699_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_1157_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1700_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .A2(_1143_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1701_ (.A1(_1154_),
    .A2(_1159_),
    .A3(_1160_),
    .B(_1161_),
    .ZN(\u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1702_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_1160_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1703_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_1147_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1704_ (.A1(_1124_),
    .A2(_1162_),
    .B(_1163_),
    .ZN(\u_arbiter.o_wb_cpu_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1705_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A4(_1157_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1706_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_1160_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1707_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .A2(_1123_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1708_ (.A1(_1154_),
    .A2(_1164_),
    .A3(_1165_),
    .B(_1166_),
    .ZN(\u_arbiter.o_wb_cpu_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1709_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_1164_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1710_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_1164_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1711_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_1123_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1712_ (.A1(_1154_),
    .A2(_1167_),
    .A3(_1168_),
    .B(_1169_),
    .ZN(\u_arbiter.o_wb_cpu_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1713_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_1167_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1714_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .A2(_1147_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1715_ (.A1(_1124_),
    .A2(_1170_),
    .B(_1171_),
    .ZN(\u_arbiter.o_wb_cpu_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1716_ (.I(_1105_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1717_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_1167_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1718_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1719_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .A2(_1147_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1720_ (.A1(_1172_),
    .A2(_1174_),
    .B(_1175_),
    .ZN(\u_arbiter.o_wb_cpu_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1721_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1722_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A4(_1164_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1723_ (.A1(_1176_),
    .A2(_1177_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1724_ (.A1(_1176_),
    .A2(_1177_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1725_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .A2(_1123_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1726_ (.A1(_1154_),
    .A2(_1178_),
    .A3(_1179_),
    .B(_1180_),
    .ZN(\u_arbiter.o_wb_cpu_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1727_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_1179_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1728_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1729_ (.A1(_1177_),
    .A2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1730_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_1123_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1731_ (.A1(_1103_),
    .A2(_1181_),
    .A3(_1183_),
    .B(_1184_),
    .ZN(\u_arbiter.o_wb_cpu_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1732_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1733_ (.A1(_1185_),
    .A2(_1183_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1734_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_1147_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1735_ (.A1(_1172_),
    .A2(_1186_),
    .B(_1187_),
    .ZN(\u_arbiter.o_wb_cpu_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1736_ (.A1(_1185_),
    .A2(_1183_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1737_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1738_ (.I(_1102_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1739_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1740_ (.A1(_1172_),
    .A2(_1189_),
    .B(_1191_),
    .ZN(\u_arbiter.o_wb_cpu_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1741_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_1185_),
    .A3(_1183_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1742_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1743_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .A2(_1190_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1744_ (.A1(_1172_),
    .A2(_1193_),
    .B(_1194_),
    .ZN(\u_arbiter.o_wb_cpu_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1745_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1746_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A4(_1183_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1747_ (.A1(_1195_),
    .A2(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1748_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_1190_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1749_ (.A1(_1172_),
    .A2(_1197_),
    .B(_1198_),
    .ZN(\u_arbiter.o_wb_cpu_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(_1195_),
    .A2(_1196_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1751_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1752_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_1190_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1753_ (.A1(_1139_),
    .A2(_1200_),
    .B(_1201_),
    .ZN(\u_arbiter.o_wb_cpu_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1754_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_1195_),
    .A3(_1196_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1755_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1756_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_1190_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1757_ (.A1(_1139_),
    .A2(_1203_),
    .B(_1204_),
    .ZN(\u_arbiter.o_wb_cpu_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1758_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A4(_1196_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1759_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1760_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_1143_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1761_ (.A1(_1139_),
    .A2(_1206_),
    .B(_1207_),
    .ZN(\u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1762_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1763_ (.A1(_1208_),
    .A2(_1205_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1764_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1765_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .I1(_1210_),
    .S(_1086_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1766_ (.I(_1211_),
    .Z(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1767_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1768_ (.I(_1212_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1769_ (.I(_1213_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1770_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1771_ (.A1(_1215_),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_1048_),
    .C(_1041_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1772_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1773_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1774_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1775_ (.A1(\u_cpu.cpu.decode.opcode[2] ),
    .A2(\u_cpu.cpu.decode.opcode[0] ),
    .A3(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1776_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1219_),
    .A3(_1220_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1777_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1220_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1778_ (.A1(\u_cpu.cpu.branch_op ),
    .A2(\u_cpu.cpu.decode.opcode[2] ),
    .A3(\u_cpu.cpu.csr_d_sel ),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1779_ (.A1(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1780_ (.A1(_1218_),
    .A2(_1221_),
    .A3(_1222_),
    .B(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1781_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1782_ (.A1(\u_cpu.rf_ram.rdata[0] ),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1783_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(\u_cpu.rf_ram_if.rtrig1 ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1784_ (.A1(\u_cpu.rf_ram_if.rtrig1 ),
    .A2(_1227_),
    .B(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1785_ (.I0(_1225_),
    .I1(_1229_),
    .S(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1786_ (.A1(_1216_),
    .A2(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1787_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1788_ (.A1(_1232_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1789_ (.A1(_1217_),
    .A2(_1231_),
    .B(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1790_ (.A1(_1214_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1791_ (.A1(_1214_),
    .A2(_1216_),
    .B(_1235_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1792_ (.I(_1045_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1793_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1794_ (.A1(_1236_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1795_ (.A1(_1236_),
    .A2(_1232_),
    .B(_1238_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1796_ (.I(_1046_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1797_ (.I(_1047_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1798_ (.A1(_1240_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1799_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1800_ (.I(_1243_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1801_ (.A1(_1244_),
    .A2(_1239_),
    .B(_1241_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1802_ (.I(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1803_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1804_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1805_ (.I(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1806_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_1053_),
    .A3(_1049_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1807_ (.A1(_1246_),
    .A2(_1247_),
    .A3(_1249_),
    .A4(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1808_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1809_ (.A1(_1218_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .B(_1248_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1810_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_1044_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1811_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(_1049_),
    .A3(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1812_ (.A1(_1213_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1813_ (.A1(_1252_),
    .A2(_1249_),
    .B(_1253_),
    .C(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1814_ (.A1(_1056_),
    .A2(_1229_),
    .B1(_1251_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1815_ (.A1(_1060_),
    .A2(_1239_),
    .A3(_1242_),
    .B1(_1245_),
    .B2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1816_ (.A1(_1078_),
    .A2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1817_ (.I(_1064_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(_1084_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1819_ (.A1(_1260_),
    .A2(_1262_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1820_ (.I(_1041_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1821_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1822_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1823_ (.A1(_1264_),
    .A2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1824_ (.A1(_1263_),
    .A2(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1825_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1826_ (.A1(_1041_),
    .A2(_1215_),
    .B1(_1268_),
    .B2(_1053_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1827_ (.A1(_1265_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1828_ (.A1(_1220_),
    .A2(_1269_),
    .A3(_1270_),
    .B(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1829_ (.I(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1830_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1831_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1832_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1833_ (.A1(_1275_),
    .A2(\u_cpu.cpu.state.init_done ),
    .A3(_1057_),
    .A4(_1042_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1834_ (.A1(_1045_),
    .A2(_1243_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1835_ (.A1(\u_cpu.cpu.branch_op ),
    .A2(_1265_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1836_ (.A1(_1060_),
    .A2(_1277_),
    .A3(_1278_),
    .B(_1264_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1837_ (.A1(_1212_),
    .A2(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1838_ (.A1(_1045_),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1839_ (.A1(_1264_),
    .A2(_1046_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1840_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_1281_),
    .A3(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1841_ (.I(\u_cpu.cpu.state.init_done ),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1842_ (.A1(_1276_),
    .A2(_1280_),
    .B1(_1283_),
    .B2(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1843_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1844_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_1286_),
    .B(_1267_),
    .C(_1225_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1845_ (.A1(_1274_),
    .A2(_1285_),
    .A3(_1267_),
    .B(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1846_ (.A1(_1273_),
    .A2(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1847_ (.I(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1848_ (.A1(_1290_),
    .A2(_1249_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1849_ (.A1(_1273_),
    .A2(_1288_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1850_ (.A1(_1289_),
    .A2(_1291_),
    .A3(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1851_ (.I(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1852_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1853_ (.A1(_1295_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .A3(_1231_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1854_ (.A1(_1049_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1855_ (.A1(_1058_),
    .A2(\u_cpu.cpu.state.init_done ),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1856_ (.A1(_1058_),
    .A2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A3(_1263_),
    .A4(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1857_ (.A1(_1212_),
    .A2(_1279_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1858_ (.A1(_1284_),
    .A2(_1283_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1859_ (.A1(_1299_),
    .A2(_1300_),
    .B(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1860_ (.A1(_1295_),
    .A2(_1230_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1861_ (.A1(_1243_),
    .A2(_1232_),
    .A3(_1230_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1862_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_1303_),
    .B(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1863_ (.A1(_1290_),
    .A2(_1248_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1864_ (.A1(_1059_),
    .A2(_1244_),
    .A3(\u_cpu.cpu.alu.cmp_r ),
    .A4(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1865_ (.A1(_1039_),
    .A2(_1302_),
    .B1(_1305_),
    .B2(_1236_),
    .C(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1866_ (.I(_1043_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1867_ (.A1(_1297_),
    .A2(_1308_),
    .B(_1309_),
    .C(_1278_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1868_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1869_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1870_ (.A1(_1311_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1871_ (.A1(_1248_),
    .A2(_1313_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1872_ (.A1(_1084_),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1873_ (.A1(_1314_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1874_ (.I(_1265_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1875_ (.A1(_1263_),
    .A2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1876_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1877_ (.A1(_1241_),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .B(\u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1878_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1879_ (.I0(_1321_),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(\u_cpu.cpu.bufreg.lsb[0] ),
    .S1(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1880_ (.A1(_1243_),
    .A2(_1320_),
    .B(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1881_ (.A1(_1243_),
    .A2(_1319_),
    .A3(_1320_),
    .B(_1323_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1882_ (.A1(_1236_),
    .A2(_1323_),
    .B(_1317_),
    .C(_1264_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1883_ (.A1(_0037_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1884_ (.A1(_1316_),
    .A2(_1318_),
    .B(_1258_),
    .C(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1885_ (.A1(_1267_),
    .A2(_1294_),
    .B(_1310_),
    .C(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1886_ (.I(_1042_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1887_ (.A1(_1274_),
    .A2(_1285_),
    .B(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1888_ (.A1(_1328_),
    .A2(_1294_),
    .B(_1329_),
    .C(_1064_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1889_ (.A1(_1064_),
    .A2(_1327_),
    .B(_1330_),
    .ZN(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1890_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1891_ (.I(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1892_ (.I(_1226_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1893_ (.A1(_1333_),
    .A2(\u_cpu.rf_ram.rdata[1] ),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1894_ (.I(_1331_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1895_ (.A1(_1335_),
    .A2(\u_cpu.rf_ram_if.rdata1[1] ),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1896_ (.A1(_1332_),
    .A2(_1334_),
    .B(_1336_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1897_ (.A1(_1333_),
    .A2(\u_cpu.rf_ram.rdata[2] ),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1898_ (.A1(_1335_),
    .A2(\u_cpu.rf_ram_if.rdata1[2] ),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1899_ (.A1(_1332_),
    .A2(_1337_),
    .B(_1338_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1900_ (.A1(_1333_),
    .A2(\u_cpu.rf_ram.rdata[3] ),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1901_ (.A1(_1335_),
    .A2(\u_cpu.rf_ram_if.rdata1[3] ),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1902_ (.A1(_1332_),
    .A2(_1339_),
    .B(_1340_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1903_ (.A1(_1226_),
    .A2(\u_cpu.rf_ram.rdata[4] ),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1904_ (.A1(_1331_),
    .A2(\u_cpu.rf_ram_if.rdata1[4] ),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1905_ (.A1(_1332_),
    .A2(_1341_),
    .B(_1342_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1906_ (.A1(_1226_),
    .A2(\u_cpu.rf_ram.rdata[5] ),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1907_ (.A1(_1331_),
    .A2(\u_cpu.rf_ram_if.rdata1[5] ),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1908_ (.A1(_1332_),
    .A2(_1343_),
    .B(_1344_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(_1226_),
    .A2(\u_cpu.rf_ram.rdata[6] ),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1910_ (.A1(_1331_),
    .A2(\u_cpu.rf_ram_if.rdata1[6] ),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1911_ (.A1(_1335_),
    .A2(_1345_),
    .B(_1346_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1912_ (.I(_1068_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1913_ (.A1(\u_cpu.rf_ram_if.rdata0[1] ),
    .A2(_1347_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1914_ (.A1(_1083_),
    .A2(_1227_),
    .B(_1348_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1915_ (.A1(\u_cpu.rf_ram_if.rdata0[2] ),
    .A2(_1347_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1916_ (.A1(_1083_),
    .A2(_1334_),
    .B(_1349_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1917_ (.I(_1067_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1918_ (.A1(\u_cpu.rf_ram_if.rdata0[3] ),
    .A2(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1919_ (.A1(_1083_),
    .A2(_1337_),
    .B(_1351_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1920_ (.A1(\u_cpu.rf_ram_if.rdata0[4] ),
    .A2(_1350_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1921_ (.A1(_1083_),
    .A2(_1339_),
    .B(_1352_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1922_ (.A1(\u_cpu.rf_ram_if.rdata0[5] ),
    .A2(_1350_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1923_ (.A1(_1347_),
    .A2(_1341_),
    .B(_1353_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1924_ (.A1(\u_cpu.rf_ram_if.rdata0[6] ),
    .A2(_1350_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1925_ (.A1(_1347_),
    .A2(_1343_),
    .B(_1354_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1926_ (.A1(\u_cpu.rf_ram_if.rdata0[7] ),
    .A2(_1350_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1927_ (.A1(_1347_),
    .A2(_1345_),
    .B(_1355_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1928_ (.I(\u_cpu.rf_ram_if.o_wen_req ),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1929_ (.A1(_1356_),
    .A2(\u_cpu.rf_ram_if.rtrig1 ),
    .A3(_1038_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1930_ (.I(_1357_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1931_ (.I0(\u_cpu.raddr[0] ),
    .I1(\u_cpu.rf_ram.i_waddr[0] ),
    .S(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1932_ (.I(_1359_),
    .Z(\u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1933_ (.I0(\u_cpu.raddr[1] ),
    .I1(\u_cpu.rf_ram.i_waddr[1] ),
    .S(_1358_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1934_ (.I(_1360_),
    .Z(\u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1935_ (.I(_1357_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1936_ (.I(_1357_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1937_ (.A1(\u_cpu.rf_ram.i_waddr[2] ),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1938_ (.A1(_1080_),
    .A2(_1361_),
    .B(_1363_),
    .ZN(\u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1939_ (.A1(\u_cpu.rf_ram.i_waddr[3] ),
    .A2(_1362_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1940_ (.A1(_1076_),
    .A2(_1361_),
    .B(_1364_),
    .ZN(\u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1941_ (.A1(\u_cpu.rf_ram.i_waddr[4] ),
    .A2(_1358_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1942_ (.A1(_1081_),
    .A2(_1361_),
    .B(_1365_),
    .ZN(\u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1943_ (.A1(\u_cpu.rf_ram.i_waddr[5] ),
    .A2(_1358_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1944_ (.A1(_1070_),
    .A2(_1361_),
    .B(_1366_),
    .ZN(\u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1945_ (.A1(\u_cpu.rf_ram.i_waddr[6] ),
    .A2(_1358_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1946_ (.A1(_1071_),
    .A2(_1362_),
    .B(_1367_),
    .ZN(\u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1947_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_1066_),
    .B1(_1362_),
    .B2(\u_cpu.rf_ram.i_waddr[7] ),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _1948_ (.I(_1368_),
    .ZN(\u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _1949_ (.I(_1361_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1950_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(_1290_),
    .A3(_1246_),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1951_ (.I(_1369_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1952_ (.A1(_1244_),
    .A2(_1040_),
    .B1(_1048_),
    .B2(_1039_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1953_ (.I(_1263_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1954_ (.I(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1955_ (.I(_1264_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1956_ (.A1(_1373_),
    .A2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1957_ (.A1(_1284_),
    .A2(_1370_),
    .A3(_1371_),
    .A4(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1958_ (.A1(_1106_),
    .A2(_1376_),
    .ZN(\u_arbiter.o_wb_cpu_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1959_ (.I(_1215_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1960_ (.A1(_1377_),
    .A2(_1087_),
    .ZN(\u_arbiter.o_wb_cpu_we ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1961_ (.I(_1302_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1962_ (.I(\u_cpu.cpu.bufreg.c_r ),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1963_ (.I(\u_cpu.cpu.decode.opcode[1] ),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1964_ (.A1(_1263_),
    .A2(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1965_ (.A1(_1328_),
    .A2(_1265_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1966_ (.A1(_1232_),
    .A2(_1381_),
    .A3(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1967_ (.A1(_1379_),
    .A2(_1383_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1968_ (.A1(_1317_),
    .A2(_1380_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1969_ (.A1(_1385_),
    .A2(_1270_),
    .B(_1306_),
    .C(_1372_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1970_ (.A1(_1309_),
    .A2(_1225_),
    .A3(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1971_ (.A1(_1384_),
    .A2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1972_ (.A1(_1379_),
    .A2(_1383_),
    .B(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1973_ (.A1(_1378_),
    .A2(_1389_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1974_ (.I(_1390_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1975_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1272_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1976_ (.A1(_1298_),
    .A2(_1279_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1977_ (.A1(_1213_),
    .A2(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1978_ (.A1(_1391_),
    .A2(_1292_),
    .B(_1393_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1979_ (.A1(_1084_),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1980_ (.A1(_1314_),
    .A2(_1315_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1981_ (.A1(_1394_),
    .A2(_1395_),
    .B(_1393_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1982_ (.I(_1370_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1983_ (.A1(_1065_),
    .A2(_1396_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1984_ (.I(_1078_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1985_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A3(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1986_ (.A1(_1317_),
    .A2(_1215_),
    .B(_1318_),
    .C(_1309_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1987_ (.I(_1392_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1988_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_1398_),
    .B(_1399_),
    .C(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1989_ (.A1(_1397_),
    .A2(_1401_),
    .B(_1396_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1990_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_1039_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1991_ (.A1(_1040_),
    .A2(_1402_),
    .B(_1240_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1992_ (.I(_1040_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1993_ (.A1(_1039_),
    .A2(_0224_),
    .B(_1240_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1994_ (.A1(_0224_),
    .A2(_1402_),
    .B(_1240_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1995_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1996_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1997_ (.I(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1998_ (.I(_0227_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1999_ (.A1(net8),
    .A2(_1086_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2000_ (.A1(_0228_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2001_ (.I(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2002_ (.A1(_1077_),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2003_ (.A1(_1298_),
    .A2(_1279_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2004_ (.A1(_1282_),
    .A2(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2005_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A4(net35),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2006_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2007_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0236_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2008_ (.A1(_0234_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2009_ (.A1(_1218_),
    .A2(_1392_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2010_ (.A1(_1282_),
    .A2(_0239_),
    .B(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2011_ (.A1(_0238_),
    .A2(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2012_ (.A1(_1059_),
    .A2(_1244_),
    .A3(_0241_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2013_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_1101_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2014_ (.A1(_1309_),
    .A2(_0242_),
    .B(_0243_),
    .C(_1328_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2015_ (.A1(_1284_),
    .A2(_1057_),
    .A3(_1369_),
    .A4(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2016_ (.A1(_0232_),
    .A2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2017_ (.A1(_0225_),
    .A2(_0246_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2018_ (.A1(_0225_),
    .A2(\u_cpu.rf_ram_if.rcnt[2] ),
    .A3(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2019_ (.A1(_0225_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2020_ (.A1(_0246_),
    .A2(_0247_),
    .A3(_0248_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2021_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0247_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2022_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0247_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2023_ (.A1(_0232_),
    .A2(_0245_),
    .A3(_0249_),
    .A4(_0250_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2024_ (.I(_0251_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2025_ (.A1(\u_cpu.raddr[1] ),
    .A2(_0249_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2026_ (.A1(_0246_),
    .A2(_0252_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2027_ (.I(\u_cpu.rf_ram.i_waddr[7] ),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2028_ (.A1(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .A2(\u_cpu.rf_ram_if.wen1_r ),
    .B1(_1038_),
    .B2(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2029_ (.I(_0254_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2030_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2031_ (.A1(_0256_),
    .A2(\u_cpu.rf_ram_if.wen0_r ),
    .A3(\u_cpu.rf_ram_if.rtrig0 ),
    .A4(_1078_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2032_ (.A1(_0253_),
    .A2(_0255_),
    .B(_0257_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2033_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0248_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2034_ (.I(_0254_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2035_ (.A1(\u_cpu.rf_ram.i_waddr[0] ),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2036_ (.A1(_0255_),
    .A2(_0258_),
    .B(_0260_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2037_ (.A1(_0225_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.raddr[0] ),
    .C(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2038_ (.A1(\u_cpu.raddr[1] ),
    .A2(_0261_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2039_ (.I(_0254_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2040_ (.I0(_0262_),
    .I1(\u_cpu.rf_ram.i_waddr[1] ),
    .S(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2041_ (.I(_0264_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2042_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2043_ (.A1(_1052_),
    .A2(_1261_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2044_ (.A1(_0265_),
    .A2(\u_cpu.cpu.immdec.imm11_7[0] ),
    .A3(_1261_),
    .B(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2045_ (.A1(\u_cpu.rf_ram.i_waddr[2] ),
    .A2(_0263_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2046_ (.A1(_0255_),
    .A2(_0267_),
    .B(_0268_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2047_ (.I(\u_cpu.rf_ram.i_waddr[3] ),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2048_ (.A1(_0256_),
    .A2(_1051_),
    .A3(_1268_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2049_ (.A1(_0256_),
    .A2(\u_cpu.cpu.immdec.imm11_7[1] ),
    .B(_0254_),
    .C(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2050_ (.A1(_0269_),
    .A2(_0255_),
    .B1(_0271_),
    .B2(_1397_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2051_ (.I(net2),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2052_ (.I(_1218_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2053_ (.A1(_0273_),
    .A2(_0233_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2054_ (.A1(_0272_),
    .A2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2055_ (.I(_0275_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2056_ (.A1(_1246_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2057_ (.A1(_1246_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2058_ (.A1(_0272_),
    .A2(_0276_),
    .A3(_0277_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2059_ (.I(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2060_ (.I(_1085_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2061_ (.A1(_0278_),
    .A2(_0277_),
    .B(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2062_ (.A1(_0278_),
    .A2(_0277_),
    .B(_0280_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2063_ (.I(_0272_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2064_ (.I(\u_cpu.cpu.mem_bytecnt[1] ),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2065_ (.A1(_0278_),
    .A2(_0277_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2066_ (.A1(_0282_),
    .A2(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2067_ (.A1(_0281_),
    .A2(_0284_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2068_ (.A1(_0272_),
    .A2(_0273_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2069_ (.I(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2070_ (.A1(_1246_),
    .A2(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2071_ (.I(\u_cpu.rf_ram_if.rgnt ),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2072_ (.A1(_0288_),
    .A2(_0245_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2073_ (.A1(_0279_),
    .A2(_1396_),
    .A3(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2074_ (.A1(_0287_),
    .A2(_0290_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2075_ (.A1(_0279_),
    .A2(_1290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2076_ (.I(_0291_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2077_ (.A1(_0281_),
    .A2(_1311_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2078_ (.A1(_1085_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2079_ (.I(_0292_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2080_ (.A1(_1077_),
    .A2(_0286_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2081_ (.A1(_1373_),
    .A2(_1374_),
    .A3(_1371_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2082_ (.A1(_0028_),
    .A2(_0294_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2083_ (.A1(_0293_),
    .A2(_0295_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2084_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_0286_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2085_ (.I(_1317_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2086_ (.A1(_1242_),
    .A2(_1277_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2087_ (.A1(_1232_),
    .A2(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2088_ (.A1(_1230_),
    .A2(_0298_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2089_ (.A1(_1234_),
    .A2(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2090_ (.A1(_0299_),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2091_ (.A1(_1236_),
    .A2(_1244_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2092_ (.A1(_0299_),
    .A2(_0301_),
    .B(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2093_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_1306_),
    .B(_0303_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2094_ (.A1(_1296_),
    .A2(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2095_ (.A1(_0302_),
    .A2(_0304_),
    .B(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2096_ (.A1(_1241_),
    .A2(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2097_ (.A1(_0297_),
    .A2(_0308_),
    .B(_0028_),
    .C(_1373_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2098_ (.A1(_0296_),
    .A2(_0309_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2099_ (.A1(_0282_),
    .A2(_1286_),
    .A3(_0035_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2100_ (.I(_0310_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2101_ (.A1(_1284_),
    .A2(_0286_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2102_ (.A1(_0281_),
    .A2(_0274_),
    .B(_0311_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2103_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_0282_),
    .B(_0278_),
    .C(\u_cpu.cpu.bufreg.lsb[0] ),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2104_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_0282_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2105_ (.A1(_1213_),
    .A2(_0312_),
    .A3(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2106_ (.A1(_1282_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2107_ (.I(_0315_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2108_ (.I(_0234_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(_1321_),
    .A2(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2110_ (.A1(_0316_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2111_ (.I(_0234_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2112_ (.I(_0243_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2113_ (.A1(net35),
    .A2(_0320_),
    .B(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2114_ (.A1(net8),
    .A2(_1101_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2115_ (.I(_0323_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2116_ (.A1(_0323_),
    .A2(_0315_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2117_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2118_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_0324_),
    .B1(_0326_),
    .B2(_1321_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2119_ (.A1(_0319_),
    .A2(_0322_),
    .B(_0327_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2120_ (.I(_0243_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2121_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_0317_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2122_ (.A1(_1321_),
    .A2(net35),
    .B(_0317_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2123_ (.A1(_0316_),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2124_ (.A1(net35),
    .A2(_0319_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2125_ (.A1(_0329_),
    .A2(_0331_),
    .B(_0321_),
    .C(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2126_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_0328_),
    .B(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2127_ (.I(_0334_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2128_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_0317_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2129_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_1321_),
    .A3(net35),
    .B(_0317_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2130_ (.A1(_0316_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2131_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_0331_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2132_ (.A1(_0335_),
    .A2(_0337_),
    .B(_0321_),
    .C(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2133_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_0328_),
    .B(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2134_ (.I(_0340_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2135_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2136_ (.I(_0323_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2137_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2138_ (.A1(_0320_),
    .A2(_0235_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2139_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_0320_),
    .B(_0316_),
    .C(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2140_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_0337_),
    .B(_0342_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2141_ (.A1(_0341_),
    .A2(_0343_),
    .B1(_0345_),
    .B2(_0346_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2142_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_0235_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2143_ (.A1(_0320_),
    .A2(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2144_ (.A1(_0243_),
    .A2(_0315_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2145_ (.I(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2146_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0320_),
    .B(_0348_),
    .C(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2147_ (.I(_0325_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2148_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_0343_),
    .B1(_0352_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2149_ (.A1(_0351_),
    .A2(_0353_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2150_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_0343_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2151_ (.I(_0325_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2152_ (.I(_0349_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2153_ (.I(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2154_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0241_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2155_ (.A1(_0354_),
    .A2(_0358_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2156_ (.I(_0325_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2157_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_0324_),
    .B1(_0350_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .C1(_0359_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2158_ (.I(_0360_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2159_ (.I(_0356_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2160_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2161_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_0343_),
    .B1(_0352_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2162_ (.A1(_0362_),
    .A2(_0363_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2163_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_0324_),
    .B1(_0326_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .C1(_0350_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2164_ (.I(_0364_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2165_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .A2(_0361_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2166_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_0343_),
    .B1(_0352_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2167_ (.A1(_0365_),
    .A2(_0366_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2168_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_0324_),
    .B1(_0326_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .C1(_0350_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2169_ (.I(_0367_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2170_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_0361_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2171_ (.I(_0342_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2172_ (.I(_0325_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2173_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_0369_),
    .B1(_0370_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2174_ (.A1(_0368_),
    .A2(_0371_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2175_ (.I(_0323_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2176_ (.I(_0356_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2177_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_0372_),
    .B1(_0326_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .C1(_0373_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2178_ (.I(_0374_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2179_ (.I(_0356_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2181_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_0369_),
    .B1(_0370_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2182_ (.A1(_0376_),
    .A2(_0377_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2183_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .A2(_0375_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2184_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_0369_),
    .B1(_0370_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(_0378_),
    .A2(_0379_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2186_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_0375_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2187_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_0369_),
    .B1(_0370_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2188_ (.A1(_0380_),
    .A2(_0381_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2189_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_0372_),
    .B1(_0326_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .C1(_0373_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2190_ (.I(_0382_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2191_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(_0375_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2192_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_0369_),
    .B1(_0370_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2193_ (.A1(_0383_),
    .A2(_0384_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2194_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_0375_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2195_ (.I(_0342_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2196_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_0386_),
    .B1(_0355_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2197_ (.A1(_0385_),
    .A2(_0387_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2198_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_0357_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2199_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_0386_),
    .B1(_0355_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2200_ (.A1(_0388_),
    .A2(_0389_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2201_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_0372_),
    .B1(_0359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .C1(_0373_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2202_ (.I(_0390_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2203_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .A2(_0357_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2204_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_0386_),
    .B1(_0355_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2205_ (.A1(_0391_),
    .A2(_0392_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2206_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_0372_),
    .B1(_0359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .C1(_0373_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2207_ (.I(_0393_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2208_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0357_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2209_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_0386_),
    .B1(_0355_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2210_ (.A1(_0394_),
    .A2(_0395_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2211_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0352_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2212_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_0386_),
    .B1(_0357_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2213_ (.A1(_0396_),
    .A2(_0397_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2214_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_0372_),
    .B1(_0359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .C1(_0373_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2215_ (.I(_0398_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2216_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2217_ (.A1(_1282_),
    .A2(_0243_),
    .A3(_0314_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2218_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_0328_),
    .B1(_0400_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2219_ (.A1(_0399_),
    .A2(_0361_),
    .B(_0401_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2220_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_0324_),
    .B1(_0350_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2221_ (.A1(_0399_),
    .A2(_0400_),
    .B(_0402_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2222_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_0342_),
    .B1(_0359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .C1(_0356_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2223_ (.I(_0403_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2224_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .A2(_0400_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2225_ (.A1(_0321_),
    .A2(_0316_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2226_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_0328_),
    .B1(_0405_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2227_ (.A1(_0404_),
    .A2(_0406_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2228_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2229_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_0328_),
    .B1(_0400_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2230_ (.A1(_0407_),
    .A2(_0361_),
    .B(_0408_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2231_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_0321_),
    .B1(_0405_),
    .B2(_1230_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2232_ (.A1(_0407_),
    .A2(_0352_),
    .B(_0409_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2233_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2234_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2235_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0410_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2236_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0410_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2237_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0410_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2238_ (.A1(_0411_),
    .A2(_0412_),
    .A3(_0413_),
    .A4(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2239_ (.I(_1090_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2240_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2241_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2242_ (.A1(_0415_),
    .A2(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2243_ (.I(_0226_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2244_ (.A1(_0417_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2245_ (.A1(_0420_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .B(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2246_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2247_ (.A1(_0419_),
    .A2(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2248_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0416_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2249_ (.A1(_1091_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2250_ (.A1(_0420_),
    .A2(\u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2251_ (.I(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2252_ (.A1(_0425_),
    .A2(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2253_ (.I(_0410_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2254_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2255_ (.I(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2256_ (.A1(_1091_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2257_ (.A1(_0417_),
    .A2(_0341_),
    .B(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2258_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0416_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2259_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_1090_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2260_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_0430_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2261_ (.I0(\u_arbiter.i_wb_cpu_rdt[2] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0430_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2262_ (.A1(_0436_),
    .A2(_0437_),
    .A3(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2263_ (.A1(_0434_),
    .A2(_0435_),
    .A3(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2264_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_1090_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2265_ (.A1(_0440_),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2266_ (.A1(_0432_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2267_ (.A1(_0429_),
    .A2(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2268_ (.I(_0438_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2269_ (.A1(_1090_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2270_ (.A1(_0226_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2271_ (.A1(_0447_),
    .A2(_0441_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2272_ (.A1(_1091_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2273_ (.A1(_0227_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2274_ (.A1(_0450_),
    .A2(_0427_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2275_ (.I0(\u_arbiter.i_wb_cpu_rdt[1] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_0416_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2276_ (.A1(_0425_),
    .A2(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2277_ (.A1(_0448_),
    .A2(_0451_),
    .B(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2278_ (.I(_0454_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2279_ (.A1(_0445_),
    .A2(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2280_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_0430_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2281_ (.A1(_0447_),
    .A2(_0441_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2282_ (.A1(_0457_),
    .A2(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2283_ (.A1(_0430_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2284_ (.A1(_0227_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2285_ (.A1(_0415_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2286_ (.A1(_0459_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2287_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2288_ (.I(_0431_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2289_ (.A1(_1091_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2290_ (.A1(_0227_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2291_ (.A1(_0465_),
    .A2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2292_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2293_ (.A1(_0450_),
    .A2(_0452_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2294_ (.I(_0470_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2295_ (.A1(_0464_),
    .A2(_0469_),
    .B(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2296_ (.A1(_0424_),
    .A2(_0444_),
    .B(_0456_),
    .C(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2297_ (.I(_0231_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2298_ (.I0(_0297_),
    .I1(_0473_),
    .S(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2299_ (.I(_0475_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(_0420_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2301_ (.A1(net8),
    .A2(_1086_),
    .A3(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2302_ (.I(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2303_ (.I(_0478_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2304_ (.I(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2305_ (.I(_0434_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2306_ (.I(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2307_ (.I(_0454_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2308_ (.I(_0483_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2309_ (.A1(_0482_),
    .A2(_0484_),
    .B1(_0469_),
    .B2(_0471_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2310_ (.I(_0478_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2311_ (.A1(_1380_),
    .A2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2312_ (.A1(_0480_),
    .A2(_0485_),
    .B(_0487_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2313_ (.A1(_0424_),
    .A2(_0428_),
    .A3(_0442_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2314_ (.I(_0450_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2315_ (.I(_0465_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2316_ (.A1(_0489_),
    .A2(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2317_ (.I(_0425_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2318_ (.I(_0447_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2319_ (.I(_0457_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2320_ (.A1(_0493_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2321_ (.I(_0441_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2322_ (.A1(_0432_),
    .A2(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2323_ (.I(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2324_ (.A1(_0495_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2325_ (.A1(_0416_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2326_ (.A1(_0227_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2327_ (.A1(_0465_),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2328_ (.A1(_0425_),
    .A2(_0452_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2329_ (.I(_0453_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2330_ (.A1(_0502_),
    .A2(_0503_),
    .B(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2331_ (.A1(_0231_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2332_ (.A1(_0492_),
    .A2(_0499_),
    .B(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2333_ (.A1(_0491_),
    .A2(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2334_ (.I(_0478_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2335_ (.A1(_0477_),
    .A2(_0505_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2336_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2337_ (.I(_0511_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2338_ (.A1(_1374_),
    .A2(_0509_),
    .B1(_0435_),
    .B2(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2339_ (.A1(_0488_),
    .A2(_0508_),
    .B(_0513_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2340_ (.I(_0230_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2341_ (.I(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2342_ (.A1(_0425_),
    .A2(_0427_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2343_ (.I(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2344_ (.A1(_0459_),
    .A2(_0462_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2345_ (.A1(_0493_),
    .A2(_0501_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2346_ (.I(_0519_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2347_ (.A1(_0468_),
    .A2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2348_ (.A1(_0448_),
    .A2(_0457_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2349_ (.I(_0411_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2350_ (.A1(_0523_),
    .A2(_0412_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2351_ (.A1(_0522_),
    .A2(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2352_ (.A1(_0518_),
    .A2(_0521_),
    .A3(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2353_ (.I(_0489_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2354_ (.I(_0501_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2355_ (.I(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2356_ (.A1(_1092_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2357_ (.A1(_0228_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2358_ (.I(_0478_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2359_ (.A1(_0527_),
    .A2(_0529_),
    .B1(_0455_),
    .B2(_0531_),
    .C(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2360_ (.A1(_0517_),
    .A2(_0526_),
    .B(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2361_ (.A1(_1377_),
    .A2(_0515_),
    .B(_0534_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2362_ (.A1(_1092_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2363_ (.A1(_0228_),
    .A2(\u_arbiter.i_wb_cpu_rdt[6] ),
    .B(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2364_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2365_ (.I(_0230_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2366_ (.A1(_1373_),
    .A2(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2367_ (.A1(_0444_),
    .A2(_0507_),
    .B1(_0512_),
    .B2(_0537_),
    .C(_0539_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2368_ (.A1(_0471_),
    .A2(_0469_),
    .B(_0483_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2369_ (.I(_0519_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2370_ (.I(_0494_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2371_ (.I(_0437_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2372_ (.A1(_0436_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2373_ (.A1(_0524_),
    .A2(_0544_),
    .B(_0448_),
    .C(_0542_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2374_ (.A1(_0438_),
    .A2(_0464_),
    .B1(_0541_),
    .B2(_0542_),
    .C(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2375_ (.A1(_0493_),
    .A2(_0501_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2376_ (.I(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2377_ (.A1(_0450_),
    .A2(_0452_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _2378_ (.A1(_0423_),
    .A2(_0540_),
    .B1(_0546_),
    .B2(_0517_),
    .C1(_0548_),
    .C2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2379_ (.A1(_0474_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2380_ (.A1(_1241_),
    .A2(_0515_),
    .B(_0551_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2381_ (.I(_0505_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2382_ (.A1(_0422_),
    .A2(_0495_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2383_ (.I(_0522_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2384_ (.A1(_0523_),
    .A2(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2385_ (.A1(_0412_),
    .A2(_0537_),
    .B(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2386_ (.A1(_0481_),
    .A2(_0464_),
    .B(_0553_),
    .C(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2387_ (.A1(_0517_),
    .A2(_0557_),
    .B(_0491_),
    .C(_0552_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2388_ (.A1(_0542_),
    .A2(_0552_),
    .B(_0558_),
    .C(_0538_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2389_ (.A1(_1240_),
    .A2(_0515_),
    .B(_0559_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2390_ (.I(_0493_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2391_ (.A1(_0536_),
    .A2(_0531_),
    .A3(_0524_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2392_ (.A1(_0435_),
    .A2(_0464_),
    .B1(_0554_),
    .B2(_0561_),
    .C(_0553_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2393_ (.A1(_0560_),
    .A2(_0453_),
    .B1(_0562_),
    .B2(_0517_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2394_ (.A1(_0474_),
    .A2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2395_ (.A1(_1059_),
    .A2(_0515_),
    .B(_0564_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2396_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_1094_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2397_ (.A1(_0445_),
    .A2(_0467_),
    .A3(_0498_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2398_ (.A1(_0422_),
    .A2(_0518_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2399_ (.A1(_0553_),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2400_ (.A1(_0492_),
    .A2(_0566_),
    .A3(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2401_ (.I(_0477_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2402_ (.I(_0528_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2403_ (.A1(_0432_),
    .A2(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2404_ (.A1(_0424_),
    .A2(_0443_),
    .B1(_0572_),
    .B2(_0438_),
    .C(_0428_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2405_ (.I(_0451_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2406_ (.I(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2407_ (.A1(_0445_),
    .A2(_0541_),
    .B(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2408_ (.A1(_0570_),
    .A2(_0504_),
    .A3(_0573_),
    .A4(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2409_ (.A1(_0511_),
    .A2(_0565_),
    .B1(_0569_),
    .B2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2410_ (.A1(_1268_),
    .A2(_0515_),
    .B(_0578_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2411_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_0486_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2412_ (.I(_0510_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2413_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_1098_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2414_ (.I(_0452_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2415_ (.A1(_0496_),
    .A2(_0494_),
    .B(_0465_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2416_ (.A1(_0481_),
    .A2(_0583_),
    .B(_0567_),
    .C(_0489_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2417_ (.A1(_0527_),
    .A2(_0481_),
    .A3(_0572_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2418_ (.A1(_0582_),
    .A2(_0584_),
    .B(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2419_ (.I(_0503_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2420_ (.A1(_0482_),
    .A2(_0541_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2421_ (.A1(_0587_),
    .A2(_0588_),
    .B(_0506_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2422_ (.A1(_0580_),
    .A2(_0581_),
    .B1(_0586_),
    .B2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2423_ (.A1(_0579_),
    .A2(_0590_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2424_ (.I(_0538_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2425_ (.I(_1093_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2426_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2427_ (.I(_0574_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2428_ (.A1(_0567_),
    .A2(_0583_),
    .B(_0470_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2429_ (.A1(_0549_),
    .A2(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2430_ (.I(_0516_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2431_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0417_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2432_ (.A1(_0598_),
    .A2(_0463_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2433_ (.I(_0435_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2434_ (.A1(_0597_),
    .A2(_0599_),
    .B(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(_0596_),
    .A2(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2436_ (.A1(_0435_),
    .A2(_0541_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2437_ (.A1(_0436_),
    .A2(_0571_),
    .B1(_0502_),
    .B2(_0593_),
    .C(_0575_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2438_ (.A1(_0594_),
    .A2(_0602_),
    .B1(_0603_),
    .B2(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2439_ (.A1(_0570_),
    .A2(_0455_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2440_ (.A1(_0511_),
    .A2(_0593_),
    .B1(_0605_),
    .B2(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2441_ (.A1(_1247_),
    .A2(_0591_),
    .B(_0607_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2442_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_1093_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2443_ (.I(_0598_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2444_ (.A1(_0465_),
    .A2(_0496_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2445_ (.A1(_0467_),
    .A2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2446_ (.A1(_0609_),
    .A2(_0611_),
    .B(_0470_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2447_ (.I(_0462_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2448_ (.A1(_0598_),
    .A2(_0613_),
    .B(_0458_),
    .C(_0494_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2449_ (.A1(_0531_),
    .A2(_0613_),
    .B(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2450_ (.A1(_0496_),
    .A2(_0494_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2451_ (.A1(_0422_),
    .A2(_0493_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2452_ (.A1(_0417_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2453_ (.A1(_0420_),
    .A2(\u_arbiter.i_wb_cpu_rdt[10] ),
    .B(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2454_ (.A1(_0411_),
    .A2(_0619_),
    .A3(_0598_),
    .A4(_0522_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2455_ (.A1(_0616_),
    .A2(_0617_),
    .B(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2456_ (.A1(_0611_),
    .A2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2457_ (.A1(_0414_),
    .A2(_0468_),
    .B1(_0519_),
    .B2(_0437_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2458_ (.I(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2459_ (.A1(_0615_),
    .A2(_0622_),
    .A3(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2460_ (.I(_0458_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2461_ (.I(_0414_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2462_ (.A1(_0438_),
    .A2(_0626_),
    .B1(_0520_),
    .B2(_0627_),
    .C(_0428_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2463_ (.A1(_0612_),
    .A2(_0625_),
    .B1(_0628_),
    .B2(_0492_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(_0503_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _2465_ (.A1(_0560_),
    .A2(_0543_),
    .B1(_0448_),
    .B2(_0608_),
    .C1(_0548_),
    .C2(_0627_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2466_ (.A1(_0630_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2467_ (.A1(_0629_),
    .A2(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2468_ (.A1(_0580_),
    .A2(_0608_),
    .B1(_0633_),
    .B2(_0606_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2469_ (.A1(_1051_),
    .A2(_0591_),
    .B(_0634_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2470_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_0479_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2471_ (.A1(_0297_),
    .A2(_1377_),
    .A3(_1044_),
    .B(_1214_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2472_ (.A1(_0570_),
    .A2(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2474_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2475_ (.A1(_0635_),
    .A2(_0638_),
    .B(_0639_),
    .C(_0578_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2476_ (.I(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2477_ (.A1(_0640_),
    .A2(_0636_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2478_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_0636_),
    .B(_0641_),
    .C(_0486_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2479_ (.A1(_0590_),
    .A2(_0642_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2480_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2481_ (.I(_0478_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2482_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0636_),
    .B(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2483_ (.A1(_0643_),
    .A2(_0638_),
    .B1(_0645_),
    .B2(_0607_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2484_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_1093_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2485_ (.A1(_0525_),
    .A2(_0599_),
    .B(_0595_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2486_ (.A1(_0543_),
    .A2(_0596_),
    .B(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2487_ (.A1(_0619_),
    .A2(_0528_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2488_ (.A1(_0490_),
    .A2(_0646_),
    .B(_0649_),
    .C(_0548_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2489_ (.A1(_0543_),
    .A2(_0610_),
    .B(_0574_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2490_ (.A1(_0575_),
    .A2(_0648_),
    .B1(_0650_),
    .B2(_0651_),
    .C(_0483_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(_0570_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2492_ (.A1(_0484_),
    .A2(_0646_),
    .B(_0652_),
    .C(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2493_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_0474_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0638_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2495_ (.A1(_0638_),
    .A2(_0654_),
    .A3(_0655_),
    .B(_0656_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2496_ (.I(_0523_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2497_ (.A1(_0657_),
    .A2(_0469_),
    .B(_0527_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2498_ (.A1(_0537_),
    .A2(_0526_),
    .B(_0599_),
    .C(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2499_ (.I(_0502_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2500_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_0592_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2501_ (.A1(_0657_),
    .A2(_0529_),
    .B1(_0660_),
    .B2(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2502_ (.A1(_0582_),
    .A2(_0537_),
    .B1(_0587_),
    .B2(_0662_),
    .C(_0504_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2503_ (.A1(_0606_),
    .A2(_0659_),
    .A3(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2504_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0532_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2505_ (.A1(_0637_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2506_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_0637_),
    .B1(_0661_),
    .B2(_0512_),
    .C(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_0664_),
    .A2(_0667_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2508_ (.A1(_0542_),
    .A2(_0613_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2509_ (.A1(_0521_),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2510_ (.A1(_0445_),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2511_ (.A1(_0609_),
    .A2(_0616_),
    .B(_0620_),
    .C(_0567_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2512_ (.A1(_0492_),
    .A2(_0670_),
    .A3(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2513_ (.I(_0506_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2514_ (.A1(_0423_),
    .A2(_0527_),
    .B1(_0582_),
    .B2(_0491_),
    .C(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2515_ (.A1(_0672_),
    .A2(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2516_ (.A1(_1372_),
    .A2(_1374_),
    .A3(_1215_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2517_ (.A1(_0297_),
    .A2(_0676_),
    .B(_1369_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2518_ (.A1(_0538_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2519_ (.A1(_0570_),
    .A2(_0677_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2520_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .S(_1095_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2521_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0678_),
    .B1(_0679_),
    .B2(\u_cpu.cpu.immdec.imm30_25[1] ),
    .C1(_0580_),
    .C2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2522_ (.A1(_0675_),
    .A2(_0681_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2523_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_0678_),
    .B1(_0679_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2524_ (.A1(_0634_),
    .A2(_0682_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2525_ (.A1(_0482_),
    .A2(_0626_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2526_ (.A1(_0436_),
    .A2(_0499_),
    .B(_0527_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2527_ (.A1(_0668_),
    .A2(_0683_),
    .B(_0684_),
    .C(_0671_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2528_ (.I(_0418_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2529_ (.A1(_0686_),
    .A2(_0520_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2530_ (.A1(_0482_),
    .A2(_0626_),
    .B(_0428_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2531_ (.I(_0418_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2532_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_0592_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2533_ (.A1(_0689_),
    .A2(_0610_),
    .B1(_0690_),
    .B2(_0660_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2534_ (.A1(_0687_),
    .A2(_0688_),
    .B1(_0691_),
    .B2(_0587_),
    .C(_0673_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2535_ (.A1(_0685_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2536_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_0678_),
    .B1(_0679_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_0690_),
    .C2(_0580_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2537_ (.A1(_0693_),
    .A2(_0694_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2538_ (.A1(_1095_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2539_ (.A1(_0228_),
    .A2(\u_arbiter.i_wb_cpu_rdt[28] ),
    .B(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2540_ (.I(_0468_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2541_ (.A1(_0413_),
    .A2(_0697_),
    .B1(_0541_),
    .B2(_0609_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2542_ (.A1(_0600_),
    .A2(_0613_),
    .B(_0614_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2543_ (.A1(_0622_),
    .A2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2544_ (.A1(_0698_),
    .A2(_0700_),
    .B(_0612_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2545_ (.A1(_1092_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2546_ (.A1(_0228_),
    .A2(\u_arbiter.i_wb_cpu_rdt[9] ),
    .B(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2547_ (.A1(_0703_),
    .A2(_0594_),
    .A3(_0548_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2548_ (.A1(_0673_),
    .A2(_0701_),
    .A3(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2549_ (.A1(_0231_),
    .A2(_0677_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2550_ (.A1(_0532_),
    .A2(_0677_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2551_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_0706_),
    .B1(_0707_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2552_ (.A1(_0512_),
    .A2(_0696_),
    .B(_0705_),
    .C(_0708_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2553_ (.I(_0412_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2554_ (.A1(_0423_),
    .A2(_0560_),
    .B(_0611_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2555_ (.A1(_0709_),
    .A2(_0469_),
    .B(_0620_),
    .C(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2556_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .S(_0592_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2557_ (.A1(_0571_),
    .A2(_0712_),
    .B(_0649_),
    .C(_0630_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2558_ (.A1(_0612_),
    .A2(_0711_),
    .B1(_0713_),
    .B2(_0490_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2559_ (.A1(_0673_),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2560_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_0706_),
    .B1(_0707_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2561_ (.A1(_0479_),
    .A2(_0552_),
    .A3(_0712_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2562_ (.A1(_0715_),
    .A2(_0716_),
    .A3(_0717_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2563_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_1098_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2564_ (.A1(_0709_),
    .A2(_0423_),
    .B(_0561_),
    .C(_0523_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2565_ (.A1(_0523_),
    .A2(_0709_),
    .B(_0554_),
    .C(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2566_ (.A1(_0689_),
    .A2(_0697_),
    .B(_0710_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2567_ (.A1(_0720_),
    .A2(_0721_),
    .B(_0612_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2568_ (.A1(_0511_),
    .A2(_0718_),
    .B1(_0722_),
    .B2(_0514_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2569_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_0678_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2570_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2571_ (.A1(_1374_),
    .A2(_0297_),
    .B(_1380_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2572_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_1223_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2573_ (.A1(_0727_),
    .A2(_0726_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2574_ (.A1(_0725_),
    .A2(_0726_),
    .B(_0728_),
    .C(_1382_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2575_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_1382_),
    .B(_0679_),
    .C(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2576_ (.A1(_0723_),
    .A2(_0724_),
    .A3(_0730_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2577_ (.A1(_0419_),
    .A2(_0609_),
    .A3(_0443_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2578_ (.A1(_0627_),
    .A2(_0442_),
    .A3(_0497_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2579_ (.A1(_0582_),
    .A2(_0731_),
    .A3(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2580_ (.A1(_1092_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2581_ (.A1(_0420_),
    .A2(\u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2582_ (.A1(_0457_),
    .A2(_0547_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2583_ (.I(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2584_ (.A1(_0609_),
    .A2(_0520_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2585_ (.A1(_0735_),
    .A2(_0432_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2586_ (.A1(_0414_),
    .A2(_0554_),
    .B1(_0739_),
    .B2(_0528_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2587_ (.A1(_0735_),
    .A2(_0737_),
    .B1(_0738_),
    .B2(_0740_),
    .C(_0597_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2588_ (.A1(_0489_),
    .A2(_0733_),
    .B(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2589_ (.A1(_0445_),
    .A2(_0571_),
    .B1(_0660_),
    .B2(_0627_),
    .C(_0575_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2590_ (.A1(_0742_),
    .A2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2591_ (.A1(_0627_),
    .A2(_0511_),
    .B1(_0744_),
    .B2(_0606_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2592_ (.A1(_1370_),
    .A2(_0727_),
    .B(_0644_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2593_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_0591_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2594_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0747_),
    .B2(_1396_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2595_ (.A1(_1309_),
    .A2(_1380_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2596_ (.A1(_1223_),
    .A2(_1266_),
    .A3(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2597_ (.A1(_1214_),
    .A2(_0749_),
    .B(_0230_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2598_ (.I(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2599_ (.I(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2600_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_0509_),
    .B(_0751_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2601_ (.A1(_0725_),
    .A2(_0752_),
    .B1(_0753_),
    .B2(_0578_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2602_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2603_ (.I(_0750_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2604_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_0509_),
    .B(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2605_ (.A1(_0754_),
    .A2(_0752_),
    .B1(_0756_),
    .B2(_0551_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2606_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2607_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_0509_),
    .B(_0755_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2608_ (.A1(_0757_),
    .A2(_0752_),
    .B1(_0758_),
    .B2(_0559_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2609_ (.I(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2610_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_0644_),
    .B(_0755_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2611_ (.A1(_0759_),
    .A2(_0752_),
    .B1(_0760_),
    .B2(_0564_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2612_ (.A1(_0703_),
    .A2(_0736_),
    .B(_0597_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2613_ (.A1(_0571_),
    .A2(_0697_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2614_ (.A1(_0598_),
    .A2(_0440_),
    .A3(_0528_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2615_ (.A1(_0549_),
    .A2(_0432_),
    .A3(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2616_ (.A1(_0761_),
    .A2(_0762_),
    .B(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2617_ (.A1(_0574_),
    .A2(_0610_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2618_ (.A1(_0553_),
    .A2(_0736_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2619_ (.A1(_0543_),
    .A2(_0464_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2620_ (.A1(_0735_),
    .A2(_0737_),
    .B1(_0767_),
    .B2(_0768_),
    .C(_0597_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2621_ (.A1(_0766_),
    .A2(_0739_),
    .B(_0769_),
    .C(_0483_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2622_ (.A1(_0735_),
    .A2(_0765_),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2623_ (.A1(_0529_),
    .A2(_0504_),
    .B(_0532_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2624_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0479_),
    .B1(_0771_),
    .B2(_0772_),
    .C(_0755_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2625_ (.A1(_1237_),
    .A2(_0752_),
    .B(_0773_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2626_ (.I(_0755_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2627_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_1093_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2628_ (.A1(_0436_),
    .A2(_0613_),
    .B(_0458_),
    .C(_0542_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2629_ (.A1(_0686_),
    .A2(_0522_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2630_ (.A1(_0687_),
    .A2(_0767_),
    .A3(_0776_),
    .A4(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2631_ (.A1(_0686_),
    .A2(_0611_),
    .B(_0778_),
    .C(_0470_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2632_ (.A1(_0549_),
    .A2(_0763_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2633_ (.A1(_0489_),
    .A2(_0490_),
    .B1(_0780_),
    .B2(_0686_),
    .C(_0503_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2634_ (.A1(_0461_),
    .A2(_0560_),
    .B(_0766_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2635_ (.A1(_0502_),
    .A2(_0775_),
    .B(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2636_ (.A1(_0779_),
    .A2(_0781_),
    .B(_0783_),
    .C(_0455_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2637_ (.A1(_0484_),
    .A2(_0775_),
    .B(_0784_),
    .C(_0653_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2638_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0514_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0774_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2640_ (.A1(_0774_),
    .A2(_0785_),
    .A3(_0786_),
    .B(_0787_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2641_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .S(_0592_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2642_ (.A1(_0413_),
    .A2(_0490_),
    .B1(_0502_),
    .B2(_0788_),
    .C(_0574_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2643_ (.A1(_0455_),
    .A2(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2644_ (.A1(_0599_),
    .A2(_0767_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2645_ (.A1(_0761_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2646_ (.A1(_0703_),
    .A2(_0765_),
    .B(_0792_),
    .C(_0594_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2647_ (.A1(_0484_),
    .A2(_0788_),
    .B1(_0790_),
    .B2(_0793_),
    .C(_0653_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2648_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0514_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2649_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0751_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2650_ (.A1(_0774_),
    .A2(_0794_),
    .A3(_0795_),
    .B(_0796_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2651_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .S(_1094_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2652_ (.A1(_0626_),
    .A2(_0697_),
    .B(_0568_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2653_ (.A1(_0619_),
    .A2(_0736_),
    .B(_0597_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2654_ (.A1(_0709_),
    .A2(_0764_),
    .B1(_0798_),
    .B2(_0799_),
    .C(_0630_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2655_ (.A1(_0560_),
    .A2(_0630_),
    .B(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2656_ (.A1(_0484_),
    .A2(_0797_),
    .B(_0801_),
    .C(_0653_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2657_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0514_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2658_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0751_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2659_ (.A1(_0774_),
    .A2(_0802_),
    .A3(_0803_),
    .B(_0804_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2660_ (.A1(_0657_),
    .A2(_0737_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2661_ (.A1(_0568_),
    .A2(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2662_ (.A1(_1094_),
    .A2(_0341_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2663_ (.A1(_1098_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_0483_),
    .C(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2664_ (.A1(_0538_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2665_ (.A1(_0657_),
    .A2(_0764_),
    .B1(_0806_),
    .B2(_0471_),
    .C(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2666_ (.A1(_1328_),
    .A2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2667_ (.A1(_0532_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2668_ (.A1(_1373_),
    .A2(_0727_),
    .B(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2669_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0751_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2670_ (.A1(_0774_),
    .A2(_0810_),
    .A3(_0813_),
    .B(_0814_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2671_ (.A1(_0553_),
    .A2(_0620_),
    .A3(_0710_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2672_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_1095_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2673_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_0509_),
    .B1(_0580_),
    .B2(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2674_ (.A1(_0480_),
    .A2(_0612_),
    .A3(_0815_),
    .B(_0817_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2675_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2676_ (.A1(_0273_),
    .A2(_1400_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2677_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2678_ (.A1(_0818_),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2679_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_1370_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2680_ (.A1(_1396_),
    .A2(_0307_),
    .B(_0821_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2681_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_1378_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2682_ (.I(_0822_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2683_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_1378_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2684_ (.I(_0823_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2685_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_1378_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2686_ (.I(_0824_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2687_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_1378_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2688_ (.I(_0825_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2689_ (.I(_1302_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2690_ (.I(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2691_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2692_ (.I(_0828_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2693_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_0827_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2694_ (.I(_0829_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2695_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_0827_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2696_ (.I(_0830_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2697_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_0827_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2698_ (.I(_0831_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2699_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_0827_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_0832_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2701_ (.I(_0826_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2702_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2703_ (.I(_0834_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2704_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_0833_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2705_ (.I(_0835_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2706_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_0833_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2707_ (.I(_0836_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2708_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_0833_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2709_ (.I(_0837_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2710_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_0833_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2711_ (.I(_0838_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2712_ (.I(_0826_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2713_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2714_ (.I(_0840_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2715_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_0839_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2716_ (.I(_0841_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2717_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_0839_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2718_ (.I(_0842_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2719_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_0839_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2720_ (.I(_0843_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2721_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_0839_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2722_ (.I(_0844_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2723_ (.I(_0826_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2724_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_0845_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2725_ (.I(_0846_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2726_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_0845_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2727_ (.I(_0847_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2728_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_0845_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2729_ (.I(_0848_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2730_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_0845_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2731_ (.I(_0849_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2732_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_0845_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2733_ (.I(_0850_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2734_ (.I(_1302_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2735_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2736_ (.I(_0852_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2737_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_0851_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2738_ (.I(_0853_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2739_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_0851_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2740_ (.I(_0854_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2741_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_0851_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2742_ (.I(_0855_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2743_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .S(_0851_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2744_ (.I(_0856_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2745_ (.A1(_1384_),
    .A2(_1387_),
    .B(_1400_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2746_ (.A1(_1384_),
    .A2(_1387_),
    .B(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2747_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_1400_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2748_ (.A1(_0826_),
    .A2(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2749_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A2(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2750_ (.A1(_1285_),
    .A2(_0858_),
    .B(_0861_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2751_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(_1290_),
    .B(_1249_),
    .C(_0233_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2752_ (.A1(_1285_),
    .A2(_0233_),
    .B(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2753_ (.A1(_1040_),
    .A2(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2754_ (.A1(_1274_),
    .A2(_0863_),
    .B(_0864_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2755_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_1400_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2756_ (.A1(_0858_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2757_ (.A1(_0863_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2758_ (.A1(_0224_),
    .A2(_0863_),
    .B(_0867_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2759_ (.A1(_1213_),
    .A2(_1392_),
    .B(net2),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2760_ (.I(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2761_ (.I(_0869_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2762_ (.A1(net2),
    .A2(_1393_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2763_ (.I(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2764_ (.I(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2765_ (.A1(_1084_),
    .A2(_0870_),
    .B1(_0873_),
    .B2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2766_ (.I(_0874_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2767_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0870_),
    .B1(_0873_),
    .B2(_1096_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2768_ (.I(_0875_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2769_ (.A1(_1096_),
    .A2(_0870_),
    .B1(_0873_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2770_ (.I(_0876_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2771_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0870_),
    .B1(_0873_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2772_ (.I(_0877_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2773_ (.I(_0869_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2774_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0878_),
    .B1(_0873_),
    .B2(_1112_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2775_ (.I(_0879_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2776_ (.I(_0872_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2777_ (.A1(_1112_),
    .A2(_0878_),
    .B1(_0880_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2778_ (.I(_0881_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2779_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_0878_),
    .B1(_0880_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2780_ (.I(_0882_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2781_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0878_),
    .B1(_0880_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2782_ (.I(_0883_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2783_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_0878_),
    .B1(_0880_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2784_ (.I(_0884_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2785_ (.I(_0868_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2786_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0885_),
    .B1(_0880_),
    .B2(_1134_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2787_ (.I(_0886_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2788_ (.I(_0872_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2789_ (.A1(_1134_),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2790_ (.I(_0888_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2791_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(_1145_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2792_ (.I(_0889_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2793_ (.A1(_1145_),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2794_ (.I(_0890_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2795_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2796_ (.I(_0891_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2797_ (.I(_0868_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2798_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0892_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2799_ (.I(_0893_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2800_ (.I(_0871_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2801_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_0892_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2802_ (.I(_0895_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2803_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0892_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2804_ (.I(_0896_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2805_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_0892_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2806_ (.I(_0897_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2807_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0892_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2808_ (.I(_0898_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2809_ (.I(_0868_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2810_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_0899_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2811_ (.I(_0900_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2812_ (.I(_0871_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2813_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2814_ (.I(_0902_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2815_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2816_ (.I(_0903_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2817_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2818_ (.I(_0904_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2819_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(_1185_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2820_ (.I(_0905_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2821_ (.I(_0868_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2822_ (.A1(_1185_),
    .A2(_0906_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2823_ (.I(_0907_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2824_ (.I(_0871_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2825_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0906_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(_0909_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2827_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0906_),
    .B1(_0908_),
    .B2(_1195_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2828_ (.I(_0910_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2829_ (.A1(_1195_),
    .A2(_0906_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2830_ (.I(_0911_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2831_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0906_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2832_ (.I(_0912_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2833_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0869_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2834_ (.I(_0913_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2835_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_0869_),
    .B1(_0872_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2836_ (.I(_0914_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2837_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_1316_),
    .B(_1050_),
    .C(_1078_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2838_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_1294_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2839_ (.A1(_1397_),
    .A2(_1050_),
    .B1(_1229_),
    .B2(_1291_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2840_ (.A1(_0916_),
    .A2(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2841_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0869_),
    .B1(_0872_),
    .B2(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2842_ (.I(_0919_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2843_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_0257_),
    .B1(_0259_),
    .B2(\u_cpu.rf_ram.i_waddr[4] ),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2844_ (.I(_0920_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2845_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0257_),
    .B1(_0259_),
    .B2(\u_cpu.rf_ram.i_waddr[5] ),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2846_ (.I(_0921_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2847_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_0257_),
    .B1(_0259_),
    .B2(\u_cpu.rf_ram.i_waddr[6] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2848_ (.I(_0922_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2849_ (.A1(_1369_),
    .A2(_1399_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2850_ (.A1(_0231_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2851_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2852_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0644_),
    .B(_0924_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2853_ (.A1(_1219_),
    .A2(_0925_),
    .B1(_0926_),
    .B2(_0745_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2854_ (.A1(_0686_),
    .A2(_0626_),
    .B1(_0520_),
    .B2(_0481_),
    .C(_0737_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2855_ (.A1(_0461_),
    .A2(_0737_),
    .B1(_0777_),
    .B2(_0927_),
    .C(_0517_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2856_ (.A1(_0630_),
    .A2(_0928_),
    .B(_0552_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2857_ (.A1(_0689_),
    .A2(_0429_),
    .A3(_0442_),
    .A4(_0498_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2858_ (.A1(_0482_),
    .A2(_0529_),
    .B1(_0660_),
    .B2(_0689_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2859_ (.A1(_0929_),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_0587_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2860_ (.A1(_0591_),
    .A2(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2861_ (.I0(\u_cpu.cpu.immdec.imm11_7[1] ),
    .I1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .S(_0923_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2862_ (.A1(_0689_),
    .A2(_0512_),
    .B1(_0934_),
    .B2(_0486_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2863_ (.A1(_0933_),
    .A2(_0935_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2864_ (.A1(_0600_),
    .A2(_0496_),
    .B1(_0498_),
    .B2(_0537_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2865_ (.A1(_0413_),
    .A2(_0660_),
    .B(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2866_ (.A1(_0413_),
    .A2(_0521_),
    .A3(_0548_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2867_ (.A1(_0603_),
    .A2(_0611_),
    .A3(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2868_ (.A1(_0761_),
    .A2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_0594_),
    .A2(_0937_),
    .B(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2870_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0479_),
    .B1(_0606_),
    .B2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2871_ (.A1(_0549_),
    .A2(_0443_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2872_ (.A1(_0454_),
    .A2(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2873_ (.A1(_0703_),
    .A2(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2874_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_0925_),
    .B1(_0945_),
    .B2(_0591_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2875_ (.A1(_0925_),
    .A2(_0942_),
    .B(_0946_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2876_ (.A1(_0582_),
    .A2(_0697_),
    .B(_0944_),
    .C(_0575_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2877_ (.A1(_0709_),
    .A2(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2878_ (.A1(_0529_),
    .A2(_0587_),
    .B1(_0554_),
    .B2(_0471_),
    .C(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2879_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_1370_),
    .A3(_1399_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2880_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0923_),
    .B(_0644_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2881_ (.A1(_0480_),
    .A2(_0949_),
    .B1(_0950_),
    .B2(_0951_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2882_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2883_ (.A1(_0492_),
    .A2(_0572_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2884_ (.A1(_0616_),
    .A2(_0953_),
    .B(_0442_),
    .C(_0594_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2885_ (.A1(_0552_),
    .A2(_0498_),
    .A3(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2886_ (.A1(_0474_),
    .A2(_0657_),
    .A3(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2887_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0486_),
    .B(_0925_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2888_ (.A1(_0952_),
    .A2(_0925_),
    .B1(_0956_),
    .B2(_0957_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2889_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_0480_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2890_ (.A1(_0723_),
    .A2(_0958_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2891_ (.A1(net8),
    .A2(\u_arbiter.o_wb_cpu_adr[1] ),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2892_ (.A1(_1095_),
    .A2(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2893_ (.A1(_0281_),
    .A2(_0960_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2894_ (.I(_0229_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2895_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2896_ (.I(_0962_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2897_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_0961_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2898_ (.I(_0963_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2899_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0961_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2900_ (.I(_0964_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2901_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_0961_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2902_ (.I(_0965_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2903_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0961_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2904_ (.I(_0966_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2905_ (.I(_0229_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2906_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2907_ (.I(_0968_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2908_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_0967_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2909_ (.I(_0969_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2910_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0967_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2911_ (.I(_0970_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2912_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_0967_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2913_ (.I(_0971_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2914_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0967_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2915_ (.I(_0972_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2916_ (.I(_0229_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2917_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2918_ (.I(_0974_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2919_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0973_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2920_ (.I(_0975_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2921_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0973_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2922_ (.I(_0976_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2923_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_0973_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2924_ (.I(_0977_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2925_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0973_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2926_ (.I(_0978_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2927_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_0229_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2928_ (.I(_0979_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2929_ (.A1(_1218_),
    .A2(_1064_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2930_ (.A1(_1214_),
    .A2(_1255_),
    .A3(_1249_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2931_ (.A1(_0980_),
    .A2(_0981_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2932_ (.I(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2933_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2934_ (.A1(_1077_),
    .A2(_0984_),
    .B(_1063_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2935_ (.A1(_0983_),
    .A2(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2936_ (.A1(_1252_),
    .A2(_0983_),
    .B(_0986_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2937_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2938_ (.A1(_1372_),
    .A2(_1377_),
    .B1(_0987_),
    .B2(_1077_),
    .C(_1063_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2939_ (.A1(_0982_),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2940_ (.A1(_0984_),
    .A2(_0983_),
    .B(_0989_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2941_ (.A1(_1275_),
    .A2(_1372_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2942_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .A2(_1397_),
    .B(_0982_),
    .C(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2943_ (.A1(_0987_),
    .A2(_0983_),
    .B(_0991_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2944_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2945_ (.A1(_1268_),
    .A2(_1062_),
    .B(_0982_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2946_ (.A1(_0992_),
    .A2(_0983_),
    .B1(_0993_),
    .B2(_1260_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2947_ (.A1(_1275_),
    .A2(_1260_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2948_ (.A1(_0273_),
    .A2(_1255_),
    .B(_1261_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2949_ (.I0(_0994_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .S(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2950_ (.I(_0996_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2951_ (.I0(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .I1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .S(_0980_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2952_ (.I(_0997_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2953_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2954_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(_0282_),
    .A3(_0278_),
    .A4(_1247_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2955_ (.A1(_1250_),
    .A2(_0277_),
    .A3(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2956_ (.A1(_1259_),
    .A2(_1000_),
    .B(_0279_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2957_ (.A1(_0998_),
    .A2(_1000_),
    .B(_1001_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2958_ (.A1(_1061_),
    .A2(_1254_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2959_ (.A1(_0273_),
    .A2(_1261_),
    .B(_1002_),
    .C(_1251_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2960_ (.A1(_1002_),
    .A2(_1259_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2961_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_1050_),
    .B(_1397_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2962_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_1003_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2963_ (.A1(_1003_),
    .A2(_1004_),
    .A3(_1005_),
    .B(_1006_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2964_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_0480_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2965_ (.A1(_0673_),
    .A2(_1007_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2966_ (.A1(_1058_),
    .A2(_0286_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2967_ (.A1(_0272_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_0820_),
    .B(_1008_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2968_ (.A1(_0653_),
    .A2(_0285_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2969_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2970_ (.A1(_0870_),
    .A2(_1009_),
    .B(_1010_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2971_ (.A1(_1333_),
    .A2(_1335_),
    .A3(\u_cpu.rf_ram.rdata[7] ),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2972_ (.I(_1011_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2973_ (.A1(_0279_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2974_ (.I(_1012_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2975_ (.A1(_0225_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2976_ (.A1(_0232_),
    .A2(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2977_ (.A1(_0245_),
    .A2(_1014_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2978_ (.A1(_1333_),
    .A2(\u_cpu.rf_ram.rdata[7] ),
    .A3(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2979_ (.I(_1015_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2980_ (.A1(_1356_),
    .A2(_1362_),
    .B(_0255_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2981_ (.A1(_0281_),
    .A2(_0232_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2982_ (.I0(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .S(_0265_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2983_ (.I0(_1016_),
    .I1(\u_cpu.rf_ram.i_wdata[0] ),
    .S(_0263_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2984_ (.I(_1017_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2985_ (.I0(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .S(_0265_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2986_ (.I0(_1018_),
    .I1(\u_cpu.rf_ram.i_wdata[1] ),
    .S(_0263_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2987_ (.I(_1019_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2988_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2989_ (.I0(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .S(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2990_ (.I(_0254_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2991_ (.I0(_1021_),
    .I1(\u_cpu.rf_ram.i_wdata[2] ),
    .S(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2992_ (.I(_1023_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2993_ (.I0(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .S(_1020_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2994_ (.I0(_1024_),
    .I1(\u_cpu.rf_ram.i_wdata[3] ),
    .S(_1022_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2995_ (.I(_1025_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2996_ (.I0(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .S(_1020_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2997_ (.I0(_1026_),
    .I1(\u_cpu.rf_ram.i_wdata[4] ),
    .S(_1022_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2998_ (.I(_1027_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2999_ (.I0(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .S(_1020_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3000_ (.I0(_1028_),
    .I1(\u_cpu.rf_ram.i_wdata[5] ),
    .S(_1022_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3001_ (.I(_1029_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3002_ (.I0(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .S(_1020_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3003_ (.I0(_1030_),
    .I1(\u_cpu.rf_ram.i_wdata[6] ),
    .S(_1022_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3004_ (.I(_1031_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3005_ (.A1(_0265_),
    .A2(\u_cpu.cpu.o_wdata0 ),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3006_ (.A1(_0256_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3007_ (.A1(\u_cpu.rf_ram.i_wdata[7] ),
    .A2(_0263_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3008_ (.A1(_0259_),
    .A2(_1032_),
    .A3(_1033_),
    .B(_1034_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3009_ (.D(_0019_),
    .CLK(net54),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3010_ (.D(_0020_),
    .CLK(net54),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3011_ (.D(_0021_),
    .CLK(net54),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3012_ (.D(_0022_),
    .CLK(net54),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3013_ (.D(_0000_),
    .CLK(net47),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3014_ (.D(_0001_),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3015_ (.D(_0002_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3016_ (.D(_0003_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3017_ (.D(_0004_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3018_ (.D(_0005_),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3019_ (.D(_0006_),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3020_ (.D(_0023_),
    .CLK(net50),
    .Q(\u_cpu.rf_ram.i_waddr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3021_ (.D(_0024_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.i_waddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3022_ (.D(_0025_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.i_waddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3023_ (.D(_0026_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.i_waddr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3024_ (.D(_0027_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.i_waddr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3025_ (.D(_0007_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3026_ (.D(_0008_),
    .CLK(net42),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3027_ (.D(_0009_),
    .CLK(net42),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3028_ (.D(_0010_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3029_ (.D(_0011_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3030_ (.D(_0012_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3031_ (.D(_0028_),
    .CLK(net72),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3032_ (.D(_0029_),
    .CLK(net76),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3033_ (.D(_0030_),
    .CLK(net74),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3034_ (.D(_0031_),
    .CLK(net74),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3035_ (.D(_0032_),
    .CLK(net76),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3036_ (.D(_0033_),
    .CLK(net76),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3037_ (.D(_0034_),
    .CLK(net76),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3038_ (.D(_0035_),
    .CLK(net74),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3039_ (.D(_0036_),
    .CLK(net72),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3040_ (.D(_0037_),
    .CLK(net74),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3041_ (.D(_0038_),
    .CLK(net72),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3042_ (.D(_0039_),
    .CLK(net75),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3043_ (.D(_0040_),
    .CLK(net73),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3044_ (.D(_0041_),
    .CLK(net86),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3045_ (.D(_0042_),
    .CLK(net86),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3046_ (.D(_0043_),
    .CLK(net114),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3047_ (.D(_0044_),
    .CLK(net86),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3048_ (.D(_0045_),
    .CLK(net87),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3049_ (.D(_0046_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3050_ (.D(_0047_),
    .CLK(net88),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3051_ (.D(_0048_),
    .CLK(net91),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3052_ (.D(_0049_),
    .CLK(net87),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3053_ (.D(_0050_),
    .CLK(net89),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3054_ (.D(_0051_),
    .CLK(net89),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3055_ (.D(_0052_),
    .CLK(net89),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3056_ (.D(_0053_),
    .CLK(net91),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3057_ (.D(_0054_),
    .CLK(net89),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3058_ (.D(_0055_),
    .CLK(net89),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3059_ (.D(_0056_),
    .CLK(net91),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3060_ (.D(_0057_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3061_ (.D(_0058_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3062_ (.D(_0059_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3063_ (.D(_0060_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3064_ (.D(_0061_),
    .CLK(net116),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3065_ (.D(_0062_),
    .CLK(net116),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3066_ (.D(_0063_),
    .CLK(net116),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3067_ (.D(_0064_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3068_ (.D(_0065_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3069_ (.D(_0066_),
    .CLK(net116),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3070_ (.D(_0067_),
    .CLK(net117),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3071_ (.D(_0068_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3072_ (.D(_0069_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3073_ (.D(_0070_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3074_ (.D(_0071_),
    .CLK(net113),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3075_ (.D(_0072_),
    .CLK(net113),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3076_ (.D(_0073_),
    .CLK(net58),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3077_ (.D(_0074_),
    .CLK(net58),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3078_ (.D(_0075_),
    .CLK(net66),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3079_ (.D(_0076_),
    .CLK(net59),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3080_ (.D(_0077_),
    .CLK(net79),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3081_ (.D(_0078_),
    .CLK(net81),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3082_ (.D(_0079_),
    .CLK(net81),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3083_ (.D(_0080_),
    .CLK(net81),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3084_ (.D(_0081_),
    .CLK(net58),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3085_ (.D(_0082_),
    .CLK(net57),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3086_ (.D(_0083_),
    .CLK(net57),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3087_ (.D(_0084_),
    .CLK(net56),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3088_ (.D(_0085_),
    .CLK(net50),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3089_ (.D(_0086_),
    .CLK(net51),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3090_ (.D(_0087_),
    .CLK(net51),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3091_ (.D(_0088_),
    .CLK(net47),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3092_ (.D(_0089_),
    .CLK(net64),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3093_ (.D(_0090_),
    .CLK(net79),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3094_ (.D(_0091_),
    .CLK(net79),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3095_ (.D(_0092_),
    .CLK(net80),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3096_ (.D(_0093_),
    .CLK(net80),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3097_ (.D(_0094_),
    .CLK(net66),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3098_ (.D(_0095_),
    .CLK(net66),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3099_ (.D(_0096_),
    .CLK(net57),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3100_ (.D(_0097_),
    .CLK(net44),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3101_ (.D(_0098_),
    .CLK(net44),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3102_ (.D(_0099_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3103_ (.D(_0100_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3104_ (.D(_0101_),
    .CLK(net49),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3105_ (.D(_0102_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3106_ (.D(_0103_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3107_ (.D(_0104_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3108_ (.D(_0105_),
    .CLK(net64),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3109_ (.D(_0106_),
    .CLK(net79),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3110_ (.D(_0107_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3111_ (.D(_0108_),
    .CLK(net73),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3112_ (.D(_0109_),
    .CLK(net100),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3113_ (.D(_0110_),
    .CLK(net100),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3114_ (.D(_0111_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3115_ (.D(_0112_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3116_ (.D(_0113_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3117_ (.D(_0114_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3118_ (.D(_0115_),
    .CLK(net76),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3119_ (.D(_0116_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3120_ (.D(_0117_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3121_ (.D(_0118_),
    .CLK(net98),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3122_ (.D(_0119_),
    .CLK(net98),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3123_ (.D(_0120_),
    .CLK(net98),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3124_ (.D(_0121_),
    .CLK(net103),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3125_ (.D(_0122_),
    .CLK(net103),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3126_ (.D(_0123_),
    .CLK(net105),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3127_ (.D(_0124_),
    .CLK(net105),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3128_ (.D(_0125_),
    .CLK(net105),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3129_ (.D(_0126_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3130_ (.D(_0127_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3131_ (.D(_0128_),
    .CLK(net108),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3132_ (.D(_0129_),
    .CLK(net108),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3133_ (.D(_0130_),
    .CLK(net108),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3134_ (.D(_0131_),
    .CLK(net108),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3135_ (.D(_0132_),
    .CLK(net108),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3136_ (.D(_0133_),
    .CLK(net119),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3137_ (.D(_0134_),
    .CLK(net119),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3138_ (.D(_0135_),
    .CLK(net118),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3139_ (.D(_0136_),
    .CLK(net118),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3140_ (.D(_0137_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3141_ (.D(_0138_),
    .CLK(net75),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3142_ (.D(_0014_),
    .CLK(net75),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3143_ (.D(_0139_),
    .CLK(net74),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3144_ (.D(_0140_),
    .CLK(net86),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3145_ (.D(_0016_),
    .CLK(net75),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3146_ (.D(_0015_),
    .CLK(net75),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3147_ (.D(_0141_),
    .CLK(net100),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3148_ (.D(_0142_),
    .CLK(net114),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3149_ (.D(_0143_),
    .CLK(net101),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3150_ (.D(_0144_),
    .CLK(net101),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3151_ (.D(_0145_),
    .CLK(net101),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3152_ (.D(_0146_),
    .CLK(net99),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3153_ (.D(_0147_),
    .CLK(net101),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3154_ (.D(_0148_),
    .CLK(net100),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3155_ (.D(_0149_),
    .CLK(net97),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3156_ (.D(_0150_),
    .CLK(net97),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3157_ (.D(_0151_),
    .CLK(net97),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3158_ (.D(_0152_),
    .CLK(net96),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3159_ (.D(_0153_),
    .CLK(net96),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3160_ (.D(_0154_),
    .CLK(net96),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3161_ (.D(_0155_),
    .CLK(net102),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3162_ (.D(_0156_),
    .CLK(net103),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3163_ (.D(_0157_),
    .CLK(net103),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3164_ (.D(_0158_),
    .CLK(net103),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3165_ (.D(_0159_),
    .CLK(net104),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3166_ (.D(_0160_),
    .CLK(net104),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3167_ (.D(_0161_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3168_ (.D(_0162_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3169_ (.D(_0163_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3170_ (.D(_0164_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3171_ (.D(_0165_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3172_ (.D(_0166_),
    .CLK(net109),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3173_ (.D(_0167_),
    .CLK(net109),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3174_ (.D(_0168_),
    .CLK(net118),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3175_ (.D(_0169_),
    .CLK(net118),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3176_ (.D(_0170_),
    .CLK(net118),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3177_ (.D(_0171_),
    .CLK(net112),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3178_ (.D(_0172_),
    .CLK(net102),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3179_ (.D(_0173_),
    .CLK(net50),
    .Q(\u_cpu.rf_ram.i_waddr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3180_ (.D(_0174_),
    .CLK(net50),
    .Q(\u_cpu.rf_ram.i_waddr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3181_ (.D(_0175_),
    .CLK(net50),
    .Q(\u_cpu.rf_ram.i_waddr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3182_ (.D(_0013_),
    .CLK(net79),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3183_ (.D(_0176_),
    .CLK(net57),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3184_ (.D(_0177_),
    .CLK(net66),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3185_ (.D(_0178_),
    .CLK(net64),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3186_ (.D(_0179_),
    .CLK(net57),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3187_ (.D(_0180_),
    .CLK(net51),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3188_ (.D(_0181_),
    .CLK(net59),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3189_ (.D(_0182_),
    .CLK(net86),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3190_ (.D(_0183_),
    .CLK(net84),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3191_ (.D(_0184_),
    .CLK(net84),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3192_ (.D(_0185_),
    .CLK(net90),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3193_ (.D(_0186_),
    .CLK(net84),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3194_ (.D(_0187_),
    .CLK(net90),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3195_ (.D(_0188_),
    .CLK(net84),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3196_ (.D(_0189_),
    .CLK(net82),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3197_ (.D(_0190_),
    .CLK(net82),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3198_ (.D(_0191_),
    .CLK(net82),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3199_ (.D(_0192_),
    .CLK(net82),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3200_ (.D(_0193_),
    .CLK(net66),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3201_ (.D(_0194_),
    .CLK(net82),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3202_ (.D(_0195_),
    .CLK(net67),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3203_ (.D(_0196_),
    .CLK(net83),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3204_ (.D(_0197_),
    .CLK(net85),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3205_ (.D(_0198_),
    .CLK(net85),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3206_ (.D(_0199_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3207_ (.D(_0200_),
    .CLK(net54),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3208_ (.D(_0201_),
    .CLK(net58),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3209_ (.D(_0202_),
    .CLK(net58),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3210_ (.D(_0203_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3211_ (.D(_0204_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3212_ (.D(_0205_),
    .CLK(net71),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3213_ (.D(_0206_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3214_ (.D(_0207_),
    .CLK(net59),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3215_ (.D(_0208_),
    .CLK(net71),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3216_ (.D(_0017_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3217_ (.D(_0209_),
    .CLK(net114),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3218_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(net36),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3219_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(net37),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3220_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(net39),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3221_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(net39),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3222_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(net39),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3223_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(net45),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3224_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(net46),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3225_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(net48),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3226_ (.D(_0210_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3227_ (.D(_0211_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3228_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(net48),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3229_ (.D(_0212_),
    .CLK(net55),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3230_ (.D(_0213_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3231_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(net36),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3232_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(net36),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3233_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(net37),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3234_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(net39),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3235_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3236_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3237_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(net45),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3238_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(net55),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3239_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(net56),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3240_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(net56),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3241_ (.D(_0214_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram_if.o_wen_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3242_ (.D(_0215_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3243_ (.D(_0216_),
    .CLK(net36),
    .Q(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3244_ (.D(_0217_),
    .CLK(net36),
    .Q(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3245_ (.D(_0218_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3246_ (.D(_0219_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3247_ (.D(_0220_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3248_ (.D(_0221_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3249_ (.D(_0222_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3250_ (.D(_0223_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__B1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__B (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__I (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__I (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__B (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__I (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__B (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__I (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A3 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__B2 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__C (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__B (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__I (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__I (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__I (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__I (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__B (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__B (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__I (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__I (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__I (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__S (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__D (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_GWEN  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[0]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[1]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[2]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[3]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[4]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[5]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[6]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[7]  (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__B (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__B (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__B (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__B (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__I0 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__B (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__B (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__B (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A3 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__B (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__S (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__S (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__S (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__S (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__S (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__B1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__B1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3410_ (.I(\u_scanchain_local.clk_out ),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3411_ (.I(\u_scanchain_local.data_out ),
    .Z(net7));
 gf180mcu_fd_ip_sram__sram256x8m8wm1 \u_cpu.rf_ram.RAM0  (.CEN(net152),
    .CLK(net44),
    .GWEN(_0018_),
    .A({\u_cpu.rf_ram.addr[7] ,
    \u_cpu.rf_ram.addr[6] ,
    \u_cpu.rf_ram.addr[5] ,
    \u_cpu.rf_ram.addr[4] ,
    \u_cpu.rf_ram.addr[3] ,
    \u_cpu.rf_ram.addr[2] ,
    \u_cpu.rf_ram.addr[1] ,
    \u_cpu.rf_ram.addr[0] }),
    .D({\u_cpu.rf_ram.i_wdata[7] ,
    \u_cpu.rf_ram.i_wdata[6] ,
    \u_cpu.rf_ram.i_wdata[5] ,
    \u_cpu.rf_ram.i_wdata[4] ,
    \u_cpu.rf_ram.i_wdata[3] ,
    \u_cpu.rf_ram.i_wdata[2] ,
    \u_cpu.rf_ram.i_wdata[1] ,
    \u_cpu.rf_ram.i_wdata[0] }),
    .Q({\u_cpu.rf_ram.rdata[7] ,
    \u_cpu.rf_ram.rdata[6] ,
    \u_cpu.rf_ram.rdata[5] ,
    \u_cpu.rf_ram.rdata[4] ,
    \u_cpu.rf_ram.rdata[3] ,
    \u_cpu.rf_ram.rdata[2] ,
    \u_cpu.rf_ram.rdata[1] ,
    \u_cpu.rf_ram.rdata[0] }),
    .WEN({_0018_,
    _0018_,
    _0018_,
    _0018_,
    _0018_,
    _0018_,
    _0018_,
    _0018_}));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.input_buf_clk  (.I(net1),
    .Z(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 \u_scanchain_local.out_flop  (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(net31),
    .Q(\u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.output_buffers[2]  (.I(\u_scanchain_local.data_out_i ),
    .Z(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.output_buffers[3]  (.I(net31),
    .Z(\u_scanchain_local.clk_out ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[0]  (.D(net3),
    .SE(net134),
    .SI(\u_arbiter.o_wb_cpu_cyc ),
    .CLK(net18),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[10]  (.D(\u_arbiter.i_wb_cpu_rdt[7] ),
    .SE(net128),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[11]  (.D(\u_arbiter.i_wb_cpu_rdt[8] ),
    .SE(net125),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(net10),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[12]  (.D(\u_arbiter.i_wb_cpu_rdt[9] ),
    .SE(net125),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[13]  (.D(\u_arbiter.i_wb_cpu_rdt[10] ),
    .SE(net128),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[14]  (.D(\u_arbiter.i_wb_cpu_rdt[11] ),
    .SE(net128),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[15]  (.D(\u_arbiter.i_wb_cpu_rdt[12] ),
    .SE(net129),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[16]  (.D(\u_arbiter.i_wb_cpu_rdt[13] ),
    .SE(net129),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[17]  (.D(\u_arbiter.i_wb_cpu_rdt[14] ),
    .SE(net129),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[18]  (.D(\u_arbiter.i_wb_cpu_rdt[15] ),
    .SE(net128),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[19]  (.D(\u_arbiter.i_wb_cpu_rdt[16] ),
    .SE(net128),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(net14),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[1]  (.D(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .SE(net134),
    .SI(\u_arbiter.o_wb_cpu_we ),
    .CLK(net18),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[20]  (.D(\u_arbiter.i_wb_cpu_rdt[17] ),
    .SE(net129),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[21]  (.D(\u_arbiter.i_wb_cpu_rdt[18] ),
    .SE(net130),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[22]  (.D(\u_arbiter.i_wb_cpu_rdt[19] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[23]  (.D(\u_arbiter.i_wb_cpu_rdt[20] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[24]  (.D(\u_arbiter.i_wb_cpu_rdt[21] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[25]  (.D(\u_arbiter.i_wb_cpu_rdt[22] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[26]  (.D(\u_arbiter.i_wb_cpu_rdt[23] ),
    .SE(net143),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(net28),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[27]  (.D(\u_arbiter.i_wb_cpu_rdt[24] ),
    .SE(net143),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(net28),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[28]  (.D(\u_arbiter.i_wb_cpu_rdt[25] ),
    .SE(net143),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(net28),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[29]  (.D(\u_arbiter.i_wb_cpu_rdt[26] ),
    .SE(net133),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[2]  (.D(net8),
    .SE(net125),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[0] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[30]  (.D(\u_arbiter.i_wb_cpu_rdt[27] ),
    .SE(net143),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(net28),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[31]  (.D(\u_arbiter.i_wb_cpu_rdt[28] ),
    .SE(net143),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(net28),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[32]  (.D(\u_arbiter.i_wb_cpu_rdt[29] ),
    .SE(net144),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(net29),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[33]  (.D(\u_arbiter.i_wb_cpu_rdt[30] ),
    .SE(net144),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(net29),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[34]  (.D(\u_arbiter.i_wb_cpu_rdt[31] ),
    .SE(net145),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[35]  (.D(\u_scanchain_local.module_data_in[34] ),
    .SE(net145),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[36]  (.D(\u_scanchain_local.module_data_in[35] ),
    .SE(net145),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[37]  (.D(\u_scanchain_local.module_data_in[36] ),
    .SE(net145),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[38]  (.D(\u_scanchain_local.module_data_in[37] ),
    .SE(net132),
    .SI(\u_arbiter.o_wb_cpu_adr[0] ),
    .CLK(net15),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[39]  (.D(\u_scanchain_local.module_data_in[38] ),
    .SE(net132),
    .SI(\u_arbiter.o_wb_cpu_adr[1] ),
    .CLK(net15),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[3]  (.D(\u_arbiter.i_wb_cpu_rdt[0] ),
    .SE(net125),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[1] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[40]  (.D(\u_scanchain_local.module_data_in[39] ),
    .SE(net145),
    .SI(\u_arbiter.o_wb_cpu_adr[2] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[41]  (.D(\u_scanchain_local.module_data_in[40] ),
    .SE(net137),
    .SI(\u_arbiter.o_wb_cpu_adr[3] ),
    .CLK(net21),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[42]  (.D(\u_scanchain_local.module_data_in[41] ),
    .SE(net137),
    .SI(\u_arbiter.o_wb_cpu_adr[4] ),
    .CLK(net21),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[43]  (.D(\u_scanchain_local.module_data_in[42] ),
    .SE(net137),
    .SI(\u_arbiter.o_wb_cpu_adr[5] ),
    .CLK(net21),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[44]  (.D(\u_scanchain_local.module_data_in[43] ),
    .SE(net138),
    .SI(\u_arbiter.o_wb_cpu_adr[6] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[45]  (.D(\u_scanchain_local.module_data_in[44] ),
    .SE(net138),
    .SI(\u_arbiter.o_wb_cpu_adr[7] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[46]  (.D(\u_scanchain_local.module_data_in[45] ),
    .SE(net135),
    .SI(\u_arbiter.o_wb_cpu_adr[8] ),
    .CLK(net20),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[47]  (.D(\u_scanchain_local.module_data_in[46] ),
    .SE(net135),
    .SI(\u_arbiter.o_wb_cpu_adr[9] ),
    .CLK(net19),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[48]  (.D(\u_scanchain_local.module_data_in[47] ),
    .SE(net135),
    .SI(\u_arbiter.o_wb_cpu_adr[10] ),
    .CLK(net19),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[49]  (.D(\u_scanchain_local.module_data_in[48] ),
    .SE(net135),
    .SI(\u_arbiter.o_wb_cpu_adr[11] ),
    .CLK(net19),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[4]  (.D(\u_arbiter.i_wb_cpu_rdt[1] ),
    .SE(net125),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[2] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[50]  (.D(\u_scanchain_local.module_data_in[49] ),
    .SE(net135),
    .SI(\u_arbiter.o_wb_cpu_adr[12] ),
    .CLK(net20),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[51]  (.D(\u_scanchain_local.module_data_in[50] ),
    .SE(net136),
    .SI(\u_arbiter.o_wb_cpu_adr[13] ),
    .CLK(net19),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[52]  (.D(\u_scanchain_local.module_data_in[51] ),
    .SE(net136),
    .SI(\u_arbiter.o_wb_cpu_adr[14] ),
    .CLK(net19),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[53]  (.D(\u_scanchain_local.module_data_in[52] ),
    .SE(net139),
    .SI(\u_arbiter.o_wb_cpu_adr[15] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[54]  (.D(\u_scanchain_local.module_data_in[53] ),
    .SE(net139),
    .SI(\u_arbiter.o_wb_cpu_adr[16] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[55]  (.D(\u_scanchain_local.module_data_in[54] ),
    .SE(net139),
    .SI(\u_arbiter.o_wb_cpu_adr[17] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[56]  (.D(\u_scanchain_local.module_data_in[55] ),
    .SE(net139),
    .SI(\u_arbiter.o_wb_cpu_adr[18] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[57]  (.D(\u_scanchain_local.module_data_in[56] ),
    .SE(net139),
    .SI(\u_arbiter.o_wb_cpu_adr[19] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[58]  (.D(\u_scanchain_local.module_data_in[57] ),
    .SE(net140),
    .SI(\u_arbiter.o_wb_cpu_adr[20] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[59]  (.D(\u_scanchain_local.module_data_in[58] ),
    .SE(net140),
    .SI(\u_arbiter.o_wb_cpu_adr[21] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[5]  (.D(\u_arbiter.i_wb_cpu_rdt[2] ),
    .SE(net126),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[3] ),
    .CLK(net10),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[60]  (.D(\u_scanchain_local.module_data_in[59] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[22] ),
    .CLK(net25),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[61]  (.D(\u_scanchain_local.module_data_in[60] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[23] ),
    .CLK(net26),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[62]  (.D(\u_scanchain_local.module_data_in[61] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[24] ),
    .CLK(net25),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[63]  (.D(\u_scanchain_local.module_data_in[62] ),
    .SE(net142),
    .SI(\u_arbiter.o_wb_cpu_adr[25] ),
    .CLK(net25),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[64]  (.D(\u_scanchain_local.module_data_in[63] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[26] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[65]  (.D(\u_scanchain_local.module_data_in[64] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[27] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[66]  (.D(\u_scanchain_local.module_data_in[65] ),
    .SE(net148),
    .SI(\u_arbiter.o_wb_cpu_adr[28] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[67]  (.D(\u_scanchain_local.module_data_in[66] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[29] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[68]  (.D(\u_scanchain_local.module_data_in[67] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[30] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[69]  (.D(\u_scanchain_local.module_data_in[68] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[31] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[6]  (.D(\u_arbiter.i_wb_cpu_rdt[3] ),
    .SE(net126),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[7]  (.D(\u_arbiter.i_wb_cpu_rdt[4] ),
    .SE(net132),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[8]  (.D(\u_arbiter.i_wb_cpu_rdt[5] ),
    .SE(net132),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[9]  (.D(\u_arbiter.i_wb_cpu_rdt[6] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout8 (.I(\u_arbiter.i_wb_cpu_ack ),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout9 (.I(net11),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout10 (.I(net11),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout11 (.I(net14),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout12 (.I(net13),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout13 (.I(net14),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout14 (.I(net17),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout15 (.I(net17),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout16 (.I(net17),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout17 (.I(net18),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout18 (.I(net34),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout19 (.I(net21),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout20 (.I(net21),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout21 (.I(net26),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout22 (.I(net26),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout23 (.I(net25),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout24 (.I(net25),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout25 (.I(net26),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout26 (.I(net33),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout27 (.I(net29),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout28 (.I(net29),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout29 (.I(net32),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout32 (.I(net33),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout33 (.I(net34),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout34 (.I(\u_scanchain_local.clk ),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout35 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout36 (.I(net38),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout38 (.I(net43),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout39 (.I(net41),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net43),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net43),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 fanout44 (.I(net69),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net53),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net53),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout48 (.I(net52),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net52),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout50 (.I(net52),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout51 (.I(net52),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout53 (.I(net62),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout54 (.I(net61),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net61),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net60),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout57 (.I(net60),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout58 (.I(net60),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net60),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net61),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net68),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net67),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net69),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout69 (.I(net124),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout70 (.I(net72),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout72 (.I(net78),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net78),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net77),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout75 (.I(net77),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net78),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net95),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout79 (.I(net81),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout81 (.I(net85),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout84 (.I(net85),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net94),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout86 (.I(net88),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net93),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout89 (.I(net91),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout90 (.I(net91),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout91 (.I(net93),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout92 (.I(net93),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout95 (.I(net123),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout96 (.I(net98),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout97 (.I(net98),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout98 (.I(net102),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout99 (.I(net100),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout100 (.I(net101),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout101 (.I(net102),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout102 (.I(net111),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net105),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net105),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net110),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net110),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout107 (.I(net109),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net110),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout110 (.I(net111),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout111 (.I(net122),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout112 (.I(net114),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout114 (.I(net117),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout115 (.I(net116),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout117 (.I(net121),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net120),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net120),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout120 (.I(net121),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout121 (.I(net122),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout122 (.I(net123),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net5),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout125 (.I(net127),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net127),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net130),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout128 (.I(net129),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net133),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout132 (.I(net133),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout133 (.I(net134),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout134 (.I(net151),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout135 (.I(net137),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout137 (.I(net142),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout138 (.I(net142),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout139 (.I(net141),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout142 (.I(net150),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout143 (.I(net146),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net146),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout145 (.I(net149),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net149),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net149),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net151),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout151 (.I(net4),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_cpu.rf_ram.RAM0_152  (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__B1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__B1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__B1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__B1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__B1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__B (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__B1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__C1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__C1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__B1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__C (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__C1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__B1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__B1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__B1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__B1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__B1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__B1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__C1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__B1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__B1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__B1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__B1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__B1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__B1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__B (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__B1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__B1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__S (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__S (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__S (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__S (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__I (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A3 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A4 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__S (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__S (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__S (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__S (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__S (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__S (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__B1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__B2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__I (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__B2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A3 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A3 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__I (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__B (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__I (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__C (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__B1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__B (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__I (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__B1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__B2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__B2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__B2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__B (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__S (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__I (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__I (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__I (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__B2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__B (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__C (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__C (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__B2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__C (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__C (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__B2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__B2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__C (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__B1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A4 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A3 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__I (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__I (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__B2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__B2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__B2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__C (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__B2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__B2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__B1 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B1 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A4 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A3 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A3 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__B (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__B2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__B (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__C (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__I (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__B2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__B2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__C (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__B1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__C (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__C (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A3 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A3 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__C (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__C1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__C1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__C2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B2 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__B (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__C (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__C (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__B (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__B1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__B (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__B1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__B1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__B (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__C (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__B (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__C (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__C (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__C (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__B (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__C (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__B (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__B1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__C2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__C1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__B2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__B2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__B1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__B2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__C (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__C (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A3 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__I (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__B (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__B (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__B1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__B2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__B2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__B2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__B2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__B (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__B (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__B (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__B (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__B (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__B (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__B2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__C2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__C (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__C (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__B (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__B (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__C (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__C (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__C (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__B1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__B1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__B2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__B1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__B1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__B2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__C (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__C (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__B (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__B1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__B1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__B2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__B2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__C1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__B1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A3 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__I (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__C (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__B2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__B (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__C (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__B (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__B (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__B1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__C (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A3 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__B2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__S (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__S (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__S (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__S (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__S (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__B1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__B1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__B2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__B (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__S (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__S (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__S (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__S (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__S (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__S (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__S (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__S (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__S (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__S (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A3 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__B2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__C (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__I (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A4 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__B1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__B (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A3 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A3 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__B (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A3 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A3 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__C (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__I (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__B (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__I (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__C (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__I (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__I (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__I (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A4 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__B (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__B2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__C (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A4 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__C (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__S (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__S (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__S (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__S (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__S (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__S (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__S (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__S (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__S (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__I (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__I (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__I (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__B (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A4 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A3 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__I (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__B (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A3 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A1 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__I (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__C (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I0 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__I (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__B1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__B2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A3 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__B2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__B (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__B (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__B (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__B (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__I (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A3 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A4 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__B (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A3 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__B (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A3 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A4 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__C (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__B (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__B2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A1 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__B (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A3 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__I (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A3 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__C (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__B (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__I (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A3 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A3 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__B1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__C (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A3 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A3 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__B2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__B (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A4 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__C (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__B (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__B (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__B2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I0 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__C (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__C (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__B (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__B (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__I (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__B1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A3 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__I (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__C (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__C (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__C (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A3 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A3 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__I (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__B2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__B (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__B (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__B2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A3 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__B (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__C (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout8_I (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__I (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__B (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__B (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__I (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__B2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_D  (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_D  (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_D  (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_D  (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_D  (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__I1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_D  (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_D  (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_D  (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_D  (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_D  (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_D  (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A2 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__A1 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_D  (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__I1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__I0 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A2 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_D  (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_D  (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_D  (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_D  (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_D  (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_D  (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_D  (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_D  (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_D  (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_D  (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_D  (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__I1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__I0 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_D  (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_D  (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_D  (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_D  (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_D  (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A2 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_D  (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_D  (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_D  (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SI  (.I(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__I (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__I (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__I (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__I (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__B (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__I (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1572__I (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__I (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A3 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_D  (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A3 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__I0 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__B2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__I0 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__I1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A3 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A2 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__I (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__B2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A2 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__D (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A2 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A2 (.I(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__B (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__I0 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[0]  (.I(\u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[1]  (.I(\u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[2]  (.I(\u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[3]  (.I(\u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[4]  (.I(\u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[5]  (.I(\u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[6]  (.I(\u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[7]  (.I(\u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__I (.I(\u_cpu.rf_ram.i_waddr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A1 (.I(\u_cpu.rf_ram.i_waddr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[0]  (.I(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__I1 (.I(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[1]  (.I(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__I1 (.I(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[2]  (.I(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__I1 (.I(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[3]  (.I(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__I1 (.I(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[4]  (.I(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__I1 (.I(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[5]  (.I(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__I1 (.I(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[6]  (.I(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__I1 (.I(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[7]  (.I(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A1 (.I(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A2 (.I(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A2 (.I(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A2 (.I(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A2 (.I(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A2 (.I(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A2 (.I(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A3 (.I(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A3 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A3 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A2 (.I(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__I (.I(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A2 (.I(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__D (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__D (.I(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__D (.I(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__D (.I(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__D (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A2 (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_D  (.I(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__B (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_D  (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_D  (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout9_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout10_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_CLK  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_CLK  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_CLK  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_CLK  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_CLK  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout12_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_CLK  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout13_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout15_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout16_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout14_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout17_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_CLK  (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_CLK  (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_CLK  (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[51]_CLK  (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[52]_CLK  (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_CLK  (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_CLK  (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_CLK  (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_CLK  (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_CLK  (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout19_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_CLK  (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_CLK  (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_CLK  (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout23_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout24_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_CLK  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_CLK  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_CLK  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_CLK  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_CLK  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_CLK  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_CLK  (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_CLK  (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout27_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.output_buffers[3]_I  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_CLKN  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout26_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_CLK  (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout77_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SE  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SE  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_SE  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_SE  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_SE  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_SE  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_SE  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SE  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_SE  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SE  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_SE  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_SE  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_SE  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_SE  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_SE  (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SE  (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_SE  (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_SE  (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_SE  (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_SE  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_SE  (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_SE  (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_SE  (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_SE  (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_SE  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_SE  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_SE  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SE  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_SE  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1758 ();
 assign io_oeb[0] = net153;
 assign io_oeb[1] = net154;
 assign io_oeb[2] = net155;
 assign io_oeb[3] = net156;
 assign io_oeb[4] = net157;
 assign io_out[2] = net158;
 assign io_out[3] = net159;
 assign io_out[4] = net160;
endmodule

