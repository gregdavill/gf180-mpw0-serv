magic
tech gf180mcuC
magscale 1 5
timestamp 1670164993
<< obsm1 >>
rect 672 1471 69328 58438
<< obsm2 >>
rect 742 569 69202 58427
<< metal3 >>
rect 69800 57792 70000 57848
rect 69800 53816 70000 53872
rect 69800 49840 70000 49896
rect 69800 45864 70000 45920
rect 69800 41888 70000 41944
rect 69800 37912 70000 37968
rect 69800 33936 70000 33992
rect 69800 29960 70000 30016
rect 69800 25984 70000 26040
rect 69800 22008 70000 22064
rect 69800 18032 70000 18088
rect 69800 14056 70000 14112
rect 69800 10080 70000 10136
rect 69800 6104 70000 6160
rect 69800 2128 70000 2184
<< obsm3 >>
rect 737 57878 69874 58422
rect 737 57762 69770 57878
rect 737 53902 69874 57762
rect 737 53786 69770 53902
rect 737 49926 69874 53786
rect 737 49810 69770 49926
rect 737 45950 69874 49810
rect 737 45834 69770 45950
rect 737 41974 69874 45834
rect 737 41858 69770 41974
rect 737 37998 69874 41858
rect 737 37882 69770 37998
rect 737 34022 69874 37882
rect 737 33906 69770 34022
rect 737 30046 69874 33906
rect 737 29930 69770 30046
rect 737 26070 69874 29930
rect 737 25954 69770 26070
rect 737 22094 69874 25954
rect 737 21978 69770 22094
rect 737 18118 69874 21978
rect 737 18002 69770 18118
rect 737 14142 69874 18002
rect 737 14026 69770 14142
rect 737 10166 69874 14026
rect 737 10050 69770 10166
rect 737 6190 69874 10050
rect 737 6074 69770 6190
rect 737 2214 69874 6074
rect 737 2098 69770 2214
rect 737 574 69874 2098
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
<< obsm4 >>
rect 4214 1508 9874 57055
rect 10094 1508 17554 57055
rect 17774 1508 25234 57055
rect 25454 1508 32914 57055
rect 33134 1508 40594 57055
rect 40814 1508 48274 57055
rect 48494 1508 55954 57055
rect 56174 1508 63634 57055
rect 63854 1508 68194 57055
rect 4214 569 68194 1508
<< labels >>
rlabel metal3 s 69800 2128 70000 2184 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 69800 6104 70000 6160 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 69800 10080 70000 10136 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 69800 14056 70000 14112 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 69800 18032 70000 18088 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 69800 41888 70000 41944 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 69800 45864 70000 45920 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 69800 49840 70000 49896 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 69800 53816 70000 53872 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 69800 57792 70000 57848 6 io_oeb[4]
port 10 nsew signal output
rlabel metal3 s 69800 22008 70000 22064 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 69800 25984 70000 26040 6 io_out[1]
port 12 nsew signal output
rlabel metal3 s 69800 29960 70000 30016 6 io_out[2]
port 13 nsew signal output
rlabel metal3 s 69800 33936 70000 33992 6 io_out[3]
port 14 nsew signal output
rlabel metal3 s 69800 37912 70000 37968 6 io_out[4]
port 15 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15129824
string GDS_FILE /home/runner/work/gf180-mpw0-serv/gf180-mpw0-serv/openlane/serv_2/runs/22_12_04_14_38/results/signoff/serv_2.magic.gds
string GDS_START 182196
<< end >>

