* NGSPICE file created from serv_2.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

.subckt serv_2 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_45_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10669__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05903_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09523__A2 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09671_ _04160_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06883_ _01452_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06337__A2 _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10023__B _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12595__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11330__A2 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08622_ _03631_ _03758_ _03763_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05834_ _01484_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08553_ u_cpu.rf_ram.memory\[54\]\[6\] _03710_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09287__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07504_ _03018_ _03015_ _03019_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08484_ _03671_ _03663_ _03672_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _02971_ _02966_ _02973_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10841__A1 u_cpu.rf_ram.memory\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09039__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07366_ _02913_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11397__A2 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__C u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09105_ _04064_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06317_ _01698_ _01962_ _01963_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07297_ _02615_ _02541_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09036_ u_cpu.rf_ram.memory\[133\]\[5\] _04019_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06248_ _01528_ _01894_ _01534_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11149__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06179_ _01600_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08014__A2 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09762__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07773__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06576__A2 _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11812__CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ _04615_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05806__I u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09869_ _02683_ _04574_ _04575_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11900_ _00422_ net89 u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12880_ _01377_ net505 u_cpu.rf_ram.memory\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11962__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11831_ _00353_ net11 u_cpu.rf_ram.memory\[68\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11543__I _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _00284_ net393 u_cpu.rf_ram.memory\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10832__A1 u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10713_ _04897_ _04711_ _04727_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12318__CLK net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11693_ _00215_ net457 u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06500__A2 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ u_cpu.rf_ram.memory\[2\]\[1\] _05185_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11388__A2 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10575_ _05143_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09450__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12314_ _00815_ net464 u_cpu.rf_ram.memory\[35\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12468__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__A2 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12245_ _00746_ net362 u_cpu.rf_ram.memory\[123\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08005__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12176_ _00690_ net425 u_cpu.rf_ram.memory\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09753__A2 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__A2 _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__A2 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11127_ _05468_ _05501_ _05503_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05870__S0 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11058_ u_cpu.rf_ram.memory\[107\]\[0\] _05458_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09505__A2 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11312__A2 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10009_ _04680_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10520__B1 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout260_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout358_I net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11076__A1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07819__A2 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout525_I net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08492__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ _02729_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ _02724_ _02728_ _02731_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08244__A2 _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06102_ _01469_ _01750_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06282__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _02678_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10051__A2 _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09992__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06033_ _01678_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11835__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10339__B1 _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11000__A1 _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07055__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09744__A2 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout105 net109 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06558__A2 _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07755__A1 u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__A2 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout127 net128 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout138 net140 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06231__B _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07984_ _03346_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09723_ _04438_ _04459_ _04466_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06935_ u_cpu.cpu.state.o_cnt_r\[1\] _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04344_ _04414_ _04421_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06866_ _02505_ u_cpu.cpu.genblk3.csr.mcause31 _02500_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07841__I _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08605_ _02943_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05817_ _01467_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09585_ u_cpu.rf_ram.memory\[121\]\[1\] _04378_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06797_ u_cpu.rf_ram.memory\[64\]\[7\] u_cpu.rf_ram.memory\[65\]\[7\] u_cpu.rf_ram.memory\[66\]\[7\]
+ u_cpu.rf_ram.memory\[67\]\[7\] _01731_ _01732_ _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11067__A1 u_cpu.rf_ram.memory\[107\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09969__S _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08536_ _03679_ _03695_ _03704_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06169__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10814__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08467_ u_cpu.rf_ram.memory\[58\]\[7\] _03649_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09680__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08483__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05916__S1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06333__I2 u_cpu.rf_ram.memory\[78\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ _02879_ _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08398_ _03568_ _03609_ _03612_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12610__CLK net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07349_ _02871_ _02893_ _02897_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09432__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06246__A1 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06192__I _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _04862_ _04963_ _05008_ _05011_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07994__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06341__S1 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ u_cpu.rf_ram.memory\[134\]\[7\] _03994_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10291_ _04925_ _04948_ _04950_ _04771_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12760__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12030_ _00544_ net420 u_cpu.rf_ram.memory\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09735__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06549__A2 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11542__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12932_ _01428_ net378 u_cpu.rf_ram.memory\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08171__A1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12863_ _01360_ net498 u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12140__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06721__A2 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__A1 u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11814_ _00336_ net16 u_cpu.rf_ram.memory\[75\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12794_ _01291_ net39 u_cpu.rf_ram.memory\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11745_ _00267_ net431 u_cpu.rf_ram.memory\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08474__A2 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09678__I _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12290__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10281__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11676_ _00198_ net466 u_cpu.rf_ram.memory\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10627_ u_cpu.rf_ram.memory\[3\]\[2\] _05176_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09423__A1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06088__I1 u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09974__A2 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10558_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _05130_ _05132_ u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout106_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10489_ _02644_ _05089_ _05090_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09726__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12228_ _00016_ net287 u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A1 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12159_ _00673_ net79 u_cpu.rf_ram.memory\[131\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10592__I0 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout475_I net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11297__A1 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06720_ u_cpu.rf_ram.memory\[128\]\[6\] u_cpu.rf_ram.memory\[129\]\[6\] u_cpu.rf_ram.memory\[130\]\[6\]
+ u_cpu.rf_ram.memory\[131\]\[6\] _01764_ _01765_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08757__I _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__A1 u_cpu.rf_ram.memory\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06651_ _02287_ _02289_ _02291_ _02293_ _01717_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06712__A2 _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11049__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09370_ _03272_ _04238_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06582_ u_cpu.rf_ram.memory\[60\]\[5\] u_cpu.rf_ram.memory\[61\]\[5\] u_cpu.rf_ram.memory\[62\]\[5\]
+ u_cpu.rf_ram.memory\[63\]\[5\] _01668_ _02034_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12633__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08321_ u_cpu.rf_ram.memory\[63\]\[7\] _03551_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08465__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06476__A1 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08252_ _03503_ _03514_ _03520_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10272__A2 _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout19_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07203_ _02721_ u_scanchain_local.module_data_in\[52\] _02722_ u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03418_ _03469_ _03475_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09414__A1 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08217__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12783__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07134_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _02716_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_dbus_dat\[14\] _02665_ _02669_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10463__S _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06016_ _01576_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12013__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06251__I1 u_cpu.rf_ram.memory\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07967_ _03333_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12163__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__A1 _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ u_cpu.rf_ram.memory\[115\]\[6\] _04451_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06918_ _02527_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07898_ _03282_ _03285_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ u_cpu.rf_ram.memory\[11\]\[6\] _04406_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06849_ _02487_ _02480_ _02488_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07900__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09568_ u_cpu.rf_ram.memory\[118\]\[2\] _04369_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _03693_ _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _04320_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__A1 u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11530_ u_cpu.rf_ram.memory\[89\]\[2\] _05758_ _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11461_ _05636_ _05707_ _05716_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08208__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10412_ _04818_ _05036_ _05045_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10015__A2 _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11392_ u_cpu.rf_ram.memory\[27\]\[3\] _05674_ _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10343_ _04683_ _04988_ _04994_ _04996_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07746__I _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09708__A2 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10274_ _04646_ _04764_ _04666_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07719__A1 u_cpu.rf_ram.memory\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12013_ _00527_ net45 u_cpu.rf_ram.memory\[141\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06078__S0 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__A1 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout480 net483 net480 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout491 net492 net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11279__A1 _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08577__I _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08144__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12915_ _01412_ net175 u_cpu.rf_ram.memory\[100\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06097__I _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12846_ _01343_ net436 u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11680__CLK net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09644__A1 u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12777_ _01274_ net12 u_cpu.rf_ram.memory\[69\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11728_ _00250_ net218 u_cpu.rf_ram.memory\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11451__A1 _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout223_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11659_ _00181_ net405 u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__A2 _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12036__CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__S1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ u_cpu.rf_ram.memory\[138\]\[1\] _03915_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08383__A1 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07821_ _03232_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07752_ u_cpu.rf_ram.memory\[41\]\[1\] _03186_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05904__I _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06703_ _01672_ _02345_ _01963_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07683_ _03139_ _03134_ _03141_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10031__B _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08686__A2 _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__S0 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ u_cpu.rf_ram.memory\[90\]\[4\] _04271_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06697__A1 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06634_ u_cpu.rf_ram.memory\[140\]\[5\] u_cpu.rf_ram.memory\[141\]\[5\] u_cpu.rf_ram.memory\[142\]\[5\]
+ u_cpu.rf_ram.memory\[143\]\[5\] _02101_ _01749_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06792__S1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09353_ _04174_ _04218_ _04226_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06565_ _02011_ _02208_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10458__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08304_ _03551_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11442__A1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09284_ u_cpu.rf_ram.memory\[123\]\[2\] _04185_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06496_ _01622_ _02140_ _01626_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06544__S1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08235_ _03349_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ u_cpu.rf_ram.memory\[6\]\[5\] _03461_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07949__A1 u_cpu.rf_ram.memory\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07117_ _02608_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12529__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08097_ u_cpu.rf_ram.memory\[74\]\[4\] _03416_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07048_ _02659_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06472__I1 u_cpu.rf_ram.memory\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11088__I _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08999_ _03735_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06775__I2 u_cpu.rf_ram.memory\[106\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10961_ _05324_ _05389_ _05396_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08677__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12700_ _01197_ net137 u_cpu.rf_ram.memory\[103\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06688__A1 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__S0 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10892_ _05350_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12631_ _01128_ net156 u_cpu.rf_ram.memory\[97\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09626__A1 u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11433__A1 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12562_ _01060_ net309 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_15_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09021__I _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11513_ _03634_ _05742_ _05748_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12493_ _00994_ net53 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06860__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11444_ _05705_ _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ _01480_ _02511_ _05664_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10326_ _04978_ _04979_ _04980_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10116__B _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10257_ _04635_ _04724_ _04703_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09691__I _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _04850_ _04853_ _04855_ _04856_ _04681_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10172__A1 _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06915__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout173_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09865__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08668__A2 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09865__B2 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06679__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12829_ _01326_ net132 u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout340_I net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09617__A1 _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout438_I net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06350_ _01985_ _01996_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09093__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06281_ u_cpu.rf_ram.memory\[48\]\[2\] u_cpu.rf_ram.memory\[49\]\[2\] u_cpu.rf_ram.memory\[50\]\[2\]
+ u_cpu.rf_ram.memory\[51\]\[2\] _01636_ _01927_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08020_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06603__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06290__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _04603_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08922_ _03932_ _03946_ _03951_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout86_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08853_ u_cpu.rf_ram.memory\[14\]\[2\] _03906_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10163__A1 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10163__B2 _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10540__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07804_ _03220_ _03212_ _03221_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12971__CLK net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ _03863_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05996_ _01499_ _01536_ _01579_ _01644_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08108__A1 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07735_ _03142_ _03170_ _03176_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09856__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08659__A2 _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07666_ u_cpu.rf_ram.memory\[46\]\[7\] _03117_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12201__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__A2 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09405_ u_cpu.rf_ram.memory\[91\]\[6\] _04254_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06617_ _01852_ _02260_ _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09608__A1 u_cpu.rf_ram.memory\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07597_ _02889_ _03081_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_94_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__A1 _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10218__A2 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09336_ _03012_ _03104_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06548_ u_cpu.rf_ram.memory\[128\]\[4\] u_cpu.rf_ram.memory\[129\]\[4\] u_cpu.rf_ram.memory\[130\]\[4\]
+ u_cpu.rf_ram.memory\[131\]\[4\] _01542_ _01760_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06517__S1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09267_ _02943_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12351__CLK net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06479_ u_cpu.rf_ram.memory\[8\]\[4\] u_cpu.rf_ram.memory\[9\]\[4\] u_cpu.rf_ram.memory\[10\]\[4\]
+ u_cpu.rf_ram.memory\[11\]\[4\] _02016_ _01507_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ _03493_ _03495_ _03497_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06842__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11919__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _04101_ _04117_ _04126_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08149_ _02889_ _02959_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07398__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11160_ u_cpu.rf_ram.memory\[84\]\[6\] _05518_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06133__C _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ _04648_ _04710_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11091_ _05211_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__A1 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04657_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10154__A1 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06453__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11993_ _00515_ net223 u_cpu.rf_ram.memory\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09847__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06205__S0 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10944_ u_cpu.rf_ram.memory\[103\]\[7\] _05375_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07322__A2 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ u_arbiter.i_wb_cpu_rdt\[27\] _05331_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11406__A1 _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12614_ _01111_ net152 u_cpu.rf_ram.memory\[93\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10209__A2 _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09075__A2 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06508__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12545_ _01045_ net254 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08822__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08590__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12476_ _00977_ net238 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12844__CLK net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11427_ u_cpu.rf_ram.memory\[25\]\[1\] _05695_ _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11358_ _05652_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10393__A1 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10309_ _04713_ _04629_ _04964_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12994__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06692__S0 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11289_ u_cpu.rf_ram.memory\[111\]\[6\] _05599_ _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A1 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13028_ _00090_ net537 u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout290_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout388_I net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06444__S0 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _01498_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12224__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09838__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07520_ _03029_ _03016_ _03030_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08765__I _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _02884_ _02957_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06402_ u_cpu.rf_ram.memory\[100\]\[3\] u_cpu.rf_ram.memory\[101\]\[3\] u_cpu.rf_ram.memory\[102\]\[3\]
+ u_cpu.rf_ram.memory\[103\]\[3\] _01934_ _01648_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ _02927_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09066__A2 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09121_ _04075_ _04065_ _04076_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06333_ u_cpu.rf_ram.memory\[76\]\[2\] u_cpu.rf_ram.memory\[77\]\[2\] u_cpu.rf_ram.memory\[78\]\[2\]
+ u_cpu.rf_ram.memory\[79\]\[2\] _01979_ _01736_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06124__I0 u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08813__A2 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06264_ u_cpu.rf_ram.memory\[32\]\[2\] u_cpu.rf_ram.memory\[33\]\[2\] u_cpu.rf_ram.memory\[34\]\[2\]
+ u_cpu.rf_ram.memory\[35\]\[2\] _01590_ _01593_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09052_ u_cpu.rf_ram.memory\[132\]\[3\] _04031_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ _03334_ _03358_ _03361_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06195_ u_cpu.rf_ram.memory\[116\]\[1\] u_cpu.rf_ram.memory\[117\]\[1\] u_cpu.rf_ram.memory\[118\]\[1\]
+ u_cpu.rf_ram.memory\[119\]\[1\] _01684_ _01685_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10384__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__S0 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _04638_ _04645_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08905_ u_cpu.rf_ram.memory\[39\]\[5\] _03933_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10136__A1 u_cpu.rf_ram.memory\[114\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09885_ _04584_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ u_cpu.rf_ram.memory\[143\]\[4\] _03893_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05938__I0 u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ _03850_ _03845_ _03852_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05979_ _01466_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09829__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ _03148_ _03156_ _03164_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08675__I _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08698_ _03730_ _03807_ _03809_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08501__A1 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07649_ _03117_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10660_ _05195_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11741__CLK net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12867__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09319_ u_cpu.rf_ram.memory\[37\]\[0\] _04206_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10591_ _05152_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10072__B1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12330_ _00831_ net454 u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12261_ _00762_ net360 u_cpu.rf_ram.memory\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08568__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ u_cpu.rf_ram.memory\[85\]\[1\] _05553_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12192_ _00706_ net268 u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput7 net7 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11143_ _02898_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07240__A1 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11074_ _05417_ _05458_ _05467_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10127__A1 _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10025_ _04713_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10678__A2 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08585__I _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11976_ _00498_ net58 u_cpu.rf_ram.memory\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09296__A2 _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10927_ _05375_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _05335_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09048__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10789_ u_cpu.rf_ram.memory\[95\]\[5\] _05287_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06806__A1 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12528_ _01029_ net324 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout303_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13022__CLK net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12459_ _00960_ net254 u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06054__B _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10366__A1 _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06665__S0 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09365__B _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout309 net312 net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_67_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07782__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__A1 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _02587_ u_cpu.rf_ram_if.rdata1\[1\] _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11614__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05902_ u_cpu.raddr\[1\] _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10090__I _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06417__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10669__A2 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _04431_ _04428_ _04432_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06882_ u_cpu.cpu.decode.opcode\[0\] _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06337__A3 _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08621_ u_cpu.rf_ram.memory\[9\]\[2\] _03762_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05833_ _01483_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06593__I0 u_cpu.rf_ram.memory\[100\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ _03675_ _03707_ _03714_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout49_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09287__A2 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11764__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05912__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07503_ u_cpu.rf_ram.memory\[20\]\[1\] _03016_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07298__A1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ u_cpu.rf_ram.memory\[57\]\[3\] _03669_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07434_ u_cpu.rf_ram.memory\[21\]\[2\] _02972_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10841__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09039__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09104_ _04063_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08798__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06316_ _01610_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07296_ _02615_ u_cpu.cpu.decode.opcode\[1\] _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09035_ _04005_ _04015_ _04022_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06247_ u_cpu.rf_ram.memory\[16\]\[2\] u_cpu.rf_ram.memory\[17\]\[2\] u_cpu.rf_ram.memory\[18\]\[2\]
+ u_cpu.rf_ram.memory\[19\]\[2\] _01529_ _01530_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07470__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06178_ _01651_ _01825_ _01654_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10357__A1 _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09211__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07222__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06656__S0 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07773__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08970__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09937_ _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09868_ u_arbiter.i_wb_cpu_rdt\[25\] _04511_ _04497_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07525__A2 _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08819_ u_cpu.rf_ram.memory\[70\]\[6\] _03880_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _04523_ _04525_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11830_ _00352_ net11 u_cpu.rf_ram.memory\[68\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _00283_ net396 u_cpu.rf_ram.memory\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _04897_ _05237_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10832__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11692_ _00214_ net456 u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ _04062_ _05184_ _05186_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _05137_ _05139_ u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12313_ _00814_ net488 u_cpu.rf_ram.memory\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07461__A1 u_cpu.rf_ram.memory\[81\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12244_ _00745_ net358 u_cpu.rf_ram.memory\[123\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10348__A1 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09202__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06647__S0 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12175_ _00689_ net424 u_cpu.rf_ram.memory\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__A1 u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11126_ u_cpu.rf_ram.memory\[69\]\[0\] _05502_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11057_ _05456_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05870__S1 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11787__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08713__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10008_ _02557_ _04677_ _04679_ _04683_ _04697_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_49_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06575__I0 u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10520__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10520__B2 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09269__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11076__A2 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout253_I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11959_ _00481_ net24 u_cpu.rf_ram.memory\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout420_I net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout518_I net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _02684_ u_scanchain_local.module_data_in\[42\] _02730_ u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09977__B1 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06101_ u_cpu.rf_ram.memory\[136\]\[0\] u_cpu.rf_ram.memory\[137\]\[0\] u_cpu.rf_ram.memory\[138\]\[0\]
+ u_cpu.rf_ram.memory\[139\]\[0\] _01747_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07081_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_dbus_dat\[21\] _02677_ _02678_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06032_ u_cpu.rf_ram.memory\[112\]\[0\] u_cpu.rf_ram.memory\[113\]\[0\] u_cpu.rf_ram.memory\[114\]\[0\]
+ u_cpu.rf_ram.memory\[115\]\[0\] _01679_ _01680_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10339__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10339__B2 _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07204__A1 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11000__A2 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12562__CLK net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06638__S0 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07394__I _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout106 net109 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout117 net122 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05907__I _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout128 net130 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout139 net140 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07983_ _02938_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09722_ u_cpu.rf_ram.memory\[116\]\[4\] _04463_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06934_ _02487_ _02571_ _02524_ _02558_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ u_cpu.rf_ram.memory\[112\]\[4\] _04418_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06865_ u_cpu.cpu.bufreg2.i_cnt_done _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10511__A1 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08604_ _03749_ _03733_ _03750_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08180__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05816_ _01466_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06810__S0 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09584_ _04332_ _04377_ _04379_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06796_ _02431_ _02433_ _02435_ _02437_ _01689_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06191__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08535_ u_cpu.rf_ram.memory\[55\]\[7\] _03693_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10814__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08466_ _03579_ _03651_ _03659_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06333__I3 u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07417_ _01463_ _02880_ _02882_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08397_ u_cpu.rf_ram.memory\[19\]\[1\] _03610_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12092__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07348_ _02892_ _02896_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10209__B _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07443__A1 u_cpu.rf_ram.memory\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\] _02827_ _02837_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07994__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ _03754_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ u_cpu.cpu.immdec.imm19_12_20\[1\] _04949_ _04947_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09196__A1 _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05817__I _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08943__A1 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10750__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12931_ _01427_ net378 u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12862_ _01359_ net496 u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06801__S0 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09024__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11813_ _00335_ net16 u_cpu.rf_ram.memory\[75\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11058__A2 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12793_ _01290_ net38 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10805__A2 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11744_ _00266_ net430 u_cpu.rf_ram.memory\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12435__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06485__A2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11675_ _00197_ net466 u_cpu.rf_ram.memory\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ _05171_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09423__A2 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__A1 u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06237__A2 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06088__I2 u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _05133_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12585__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07985__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10488_ _02635_ _05089_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12227_ _00015_ net287 u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12158_ _00672_ net78 u_cpu.rf_ram.memory\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10741__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10592__I1 _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11109_ _05473_ _05489_ _05492_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12089_ _00603_ net72 u_cpu.rf_ram.memory\[138\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout370_I net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11297__A2 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06548__I0 u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11464__I _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout468_I net469 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06650_ _02006_ _02292_ _01728_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11049__A2 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06581_ _02218_ _02220_ _02222_ _02224_ _01665_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_80_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09111__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08320_ _03509_ _03553_ _03561_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06476__A2 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08251_ u_cpu.rf_ram.memory\[65\]\[3\] _03518_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__I0 u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11802__CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07389__I _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06507__B _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07202_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _02772_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ u_cpu.rf_ram.memory\[68\]\[3\] _03473_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09414__A2 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07133_ _02715_ _02710_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ _02668_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11952__CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10980__A1 u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09178__A1 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06015_ _01660_ _01662_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__I _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__B _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09109__I _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06400__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06251__I2 u_cpu.rf_ram.memory\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07966_ _02913_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09705_ _04440_ _04448_ _04455_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06917_ _02518_ _02554_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07897_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _03284_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09350__A1 u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09636_ _04077_ _04403_ _04410_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06848_ _02487_ _01439_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12458__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09567_ _04364_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06779_ _01582_ _02420_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08518_ _03693_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04251_ _04321_ _04324_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10799__A1 _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06467__A2 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _03101_ _03595_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11460__A2 _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11460_ u_cpu.rf_ram.memory\[24\]\[7\] _05705_ _05716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09405__A2 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10411_ u_cpu.rf_ram.memory\[31\]\[7\] _05034_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11212__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11391_ _05625_ _05670_ _05675_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10342_ _04952_ _04995_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10971__A1 _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11549__I _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10273_ _04724_ _04762_ _04933_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12012_ _00526_ net61 u_cpu.rf_ram.memory\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06078__S1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10723__A1 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06778__I0 u_cpu.rf_ram.memory\[124\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__A2 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout470 net495 net470 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout481 net483 net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_65_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout492 net493 net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09341__A1 u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12914_ _01411_ net196 u_cpu.rf_ram.memory\[100\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06378__I _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__A2 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12845_ _01342_ net435 u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08593__I _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12776_ _01273_ net13 u_cpu.rf_ram.memory\[69\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11727_ _00249_ net210 u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11451__A2 _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06702__I0 u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11658_ _00180_ net404 u_cpu.rf_ram.memory\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11975__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ u_cpu.rf_ram.memory\[109\]\[3\] _05164_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout216_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11589_ _00111_ net410 u_cpu.rf_ram.memory\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__A4 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A2 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__I2 u_cpu.rf_ram.memory\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10714__A1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07820_ _03232_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09580__A1 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08383__A2 _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08768__I _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10190__A2 _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ _03129_ _03185_ _03187_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06784__I3 u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__B _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06702_ u_cpu.rf_ram.memory\[88\]\[6\] u_cpu.rf_ram.memory\[89\]\[6\] u_cpu.rf_ram.memory\[90\]\[6\]
+ u_cpu.rf_ram.memory\[91\]\[6\] _01961_ _01674_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08135__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ u_cpu.rf_ram.memory\[45\]\[2\] _03140_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09883__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09421_ _04256_ _04267_ _04273_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06633_ _02188_ _02276_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06241__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12750__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ u_cpu.rf_ram.memory\[36\]\[6\] _04221_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06564_ u_cpu.rf_ram.memory\[4\]\[5\] u_cpu.rf_ram.memory\[5\]\[5\] u_cpu.rf_ram.memory\[6\]\[5\]
+ u_cpu.rf_ram.memory\[7\]\[5\] _01782_ _01897_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09635__A2 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05920__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _03550_ _03231_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11442__A2 _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ _04180_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06495_ u_cpu.rf_ram.memory\[56\]\[4\] u_cpu.rf_ram.memory\[57\]\[4\] u_cpu.rf_ram.memory\[58\]\[4\]
+ u_cpu.rf_ram.memory\[59\]\[4\] _01623_ _01812_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ _03507_ _03496_ _03508_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08165_ _02934_ _03457_ _03464_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10474__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07949__A2 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07116_ _02698_ _02700_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08071__A1 _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ _03343_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07047_ u_arbiter.i_wb_cpu_rdt\[9\] u_arbiter.i_wb_cpu_dbus_dat\[6\] _02658_ _02659_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10705__A1 _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09571__A1 _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ _03993_ _03995_ _03997_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12280__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ u_cpu.rf_ram.memory\[17\]\[4\] _03318_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06775__I3 u_cpu.rf_ram.memory\[107\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11848__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08126__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10960_ u_cpu.rf_ram.memory\[104\]\[5\] _05392_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06527__I3 u_cpu.rf_ram.memory\[83\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09619_ _04081_ _04390_ _04399_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06688__A2 _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__S1 _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10891_ _05315_ _05351_ _05354_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12630_ _01127_ net159 u_cpu.rf_ram.memory\[97\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09626__A2 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07637__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12561_ _01059_ net309 u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11433__A2 _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11512_ u_cpu.rf_ram.memory\[100\]\[3\] _05746_ _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12492_ _00993_ net237 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11443_ _05705_ _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06860__A2 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11374_ _05657_ _01480_ _02515_ _05663_ _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _04790_ _04688_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10116__C _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10256_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _04774_ _04918_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12623__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08365__A2 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__I _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _04729_ _04821_ _04849_ _04664_ _04790_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A2 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__A2 _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12773__CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09865__A2 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07876__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__A2 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12828_ _01325_ net125 u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12003__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09617__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07628__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout333_I net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12759_ _01256_ net207 u_cpu.rf_ram.memory\[83\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06280_ _01637_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout500_I net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12153__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11188__A1 u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10935__A1 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout8 net9 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10093__I _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _04658_ _04660_ _04661_ _04607_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_89_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ u_cpu.rf_ram.memory\[137\]\[2\] _03950_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09553__A1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _03901_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10821__I _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06367__A1 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__B _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__I _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10163__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout79_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11360__B2 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07803_ u_cpu.rf_ram.memory\[48\]\[3\] _03218_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08783_ _03052_ _03395_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05995_ _01580_ _01614_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_22_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08108__A2 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ u_cpu.rf_ram.memory\[51\]\[3\] _03174_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11112__A1 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07665_ _03029_ _03119_ _03127_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10469__S _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09404_ _04173_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ u_cpu.rf_ram.memory\[80\]\[5\] u_cpu.rf_ram.memory\[81\]\[5\] u_cpu.rf_ram.memory\[82\]\[5\]
+ u_cpu.rf_ram.memory\[83\]\[5\] _01584_ _01965_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ _02879_ _02883_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09122__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07619__A1 u_cpu.rf_ram.memory\[78\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09335_ _04177_ _04206_ _04215_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11415__A2 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06547_ _01752_ _02191_ _01756_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08292__A1 u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09266_ _04171_ _04155_ _04172_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06478_ _01785_ _02122_ _01902_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08217_ u_cpu.rf_ram.memory\[66\]\[0\] _03496_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09197_ u_cpu.rf_ram.memory\[127\]\[7\] _04115_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11179__A1 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08044__A1 u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ _03426_ _03443_ _03452_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12646__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10926__A1 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06414__C _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09792__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08595__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ _03353_ _03398_ _03407_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10110_ _04721_ _04713_ _04616_ _04789_ _04777_ _04661_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_1_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11090_ _05478_ _05470_ _05479_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11670__CLK net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09544__A1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08347__A2 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12796__CLK net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _04622_ _04623_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06453__S1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11992_ _00514_ net223 u_cpu.rf_ram.memory\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11103__A1 _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12026__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10943_ _05326_ _05377_ _05385_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06205__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07322__A3 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10874_ _05344_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12613_ _01110_ net151 u_cpu.rf_ram.memory\[93\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11406__A2 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10465__I0 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12544_ _01044_ net255 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10906__I _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12475_ _00976_ net237 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06605__B _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11426_ _05618_ _05694_ _05696_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08586__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11357_ _05651_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _05640_ _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06141__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10393__A2 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10308_ _04636_ _04822_ _04624_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11288_ _05564_ _05596_ _05603_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06692__S1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__A1 u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13027_ _00089_ net529 u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08338__A2 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10641__I _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _04897_ _04902_ _04821_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06349__A1 _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10145__A2 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11342__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06444__S1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09838__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout450_I net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12519__CLK net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ _02982_ _02967_ _02983_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ _01499_ _02010_ _02021_ _02046_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_56_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _02926_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ u_cpu.rf_ram.memory\[12\]\[4\] _04071_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06332_ _01502_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08274__A1 _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__I1 u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10081__A1 _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09051_ _04000_ _04027_ _04032_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06263_ _01796_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06824__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ u_cpu.rf_ram.memory\[119\]\[1\] _03359_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06194_ _01678_ _01841_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10908__A1 u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _04644_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06683__S1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08904_ _03748_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11333__A1 u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09884_ _02984_ _04426_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ _03853_ _03889_ _03895_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05938__I1 u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ u_cpu.rf_ram.memory\[73\]\[2\] _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05978_ _01622_ _01625_ _01626_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09829__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ u_cpu.rf_ram.memory\[44\]\[6\] _03159_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12199__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ u_cpu.rf_ram.memory\[140\]\[0\] _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08501__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ _03083_ _03104_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07579_ u_cpu.rf_ram.memory\[80\]\[0\] _03071_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _04204_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08265__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10590_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _05107_ _05110_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10072__A1 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09249_ _04158_ _04154_ _04159_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06371__S0 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06425__B _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08017__A1 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12260_ _00761_ net355 u_cpu.rf_ram.memory\[37\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11211_ _05201_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12191_ _00705_ net260 u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11572__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11142_ _05486_ _05502_ _05511_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06674__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11073_ u_cpu.rf_ram.memory\[107\]\[7\] _05456_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11324__A1 u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10127__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10024_ _04630_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11975_ _00497_ net31 u_cpu.rf_ram.memory\[52\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10926_ _03052_ _05374_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10857_ _05330_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09697__I _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10788_ _05212_ _05283_ _05290_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12527_ _01028_ net324 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout129_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12961__CLK net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08008__A1 _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12458_ _00959_ net253 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11409_ _05681_ _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12389_ _00890_ net474 u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06665__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout498_I net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ _02583_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10118__A2 _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05901_ _01549_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06881_ _02517_ _02514_ _02519_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06417__S1 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _03757_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12341__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08731__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05832_ _01477_ _01482_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07680__I _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11909__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08551_ u_cpu.rf_ram.memory\[54\]\[5\] _03710_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10320__B _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07502_ _02914_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08482_ _03340_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12491__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07433_ _02965_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08247__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07364_ _02902_ u_cpu.rf_ram_if.wdata0_r\[1\] _02911_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_50_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09103_ _03256_ _03153_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout8_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06315_ u_cpu.rf_ram.memory\[88\]\[2\] u_cpu.rf_ram.memory\[89\]\[2\] u_cpu.rf_ram.memory\[90\]\[2\]
+ u_cpu.rf_ram.memory\[91\]\[2\] _01961_ _01700_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09995__A1 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08798__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ _02763_ _02848_ _02849_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09034_ u_cpu.rf_ram.memory\[133\]\[4\] _04019_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06246_ _01890_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09747__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06177_ u_cpu.rf_ram.memory\[96\]\[1\] u_cpu.rf_ram.memory\[97\]\[1\] u_cpu.rf_ram.memory\[98\]\[1\]
+ u_cpu.rf_ram.memory\[99\]\[1\] _01652_ _01824_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11554__A1 u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10357__A2 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06656__S1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08970__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ _04613_ _04627_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11306__A1 _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__A1 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09867_ _04491_ _04486_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08818_ _03857_ _03877_ _03884_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11589__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09798_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _04497_ _04524_ _03289_ _04525_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12834__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ u_cpu.rf_ram.memory\[72\]\[5\] _03836_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11760_ _00282_ net396 u_cpu.rf_ram.memory\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10711_ _04728_ _04666_ _04739_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ _00213_ net456 u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10642_ u_cpu.rf_ram.memory\[2\]\[0\] _05185_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10573_ _05142_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12312_ _00813_ net488 u_cpu.rf_ram.memory\[35\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07461__A2 _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12243_ _00744_ net358 u_cpu.rf_ram.memory\[123\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10348__A2 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12174_ _00688_ net424 u_cpu.rf_ram.memory\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08410__A1 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06647__S1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11125_ _05500_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08961__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11056_ _05456_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10007_ _04685_ _04688_ _04696_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08713__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10520__A2 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08477__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11958_ _00480_ net24 u_cpu.rf_ram.memory\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07005__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10284__A1 _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10909_ _05309_ _05363_ _05365_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout246_I net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11889_ _00411_ net270 u_cpu.rf_ram.memory\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10036__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09977__A1 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout413_I net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09977__B2 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06100_ _01748_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_12_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ _02664_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06031_ _01585_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09729__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12707__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11536__A1 u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10339__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08401__A1 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06638__S1 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__C _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout107 net109 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net120 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout129 net130 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07982_ _03344_ _03330_ _03345_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _04436_ _04459_ _04465_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06933_ _02568_ _02569_ _02571_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12857__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09901__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08704__A2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06864_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _04342_ _04414_ _04420_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05923__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05815_ _01439_ _01440_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08603_ u_cpu.rf_ram.memory\[52\]\[5\] _03740_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09583_ u_cpu.rf_ram.memory\[121\]\[0\] _04378_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06795_ _02082_ _02436_ _02085_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__S1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06191__A2 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11881__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _03677_ _03695_ _03703_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08468__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ u_cpu.rf_ram.memory\[58\]\[6\] _03654_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07416_ _02888_ _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12237__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ _03563_ _03609_ _03611_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07691__A2 _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07347_ _02894_ _02895_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__S0 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08640__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07278_ _02832_ _02827_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _04009_ _03996_ _04010_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06229_ _01469_ _01876_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11527__A1 u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09196__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__B _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08943__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06954__A1 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__A2 _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ _02706_ _02642_ _04610_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12930_ _01426_ net378 u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10502__A2 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05833__I _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12861_ _01358_ net317 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06801__S1 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13012__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11812_ _00334_ net34 u_cpu.rf_ram.memory\[75\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08459__A1 u_cpu.rf_ram.memory\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12792_ _01289_ net70 u_cpu.rf_ram.memory\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09120__A2 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11743_ _00265_ net430 u_cpu.rf_ram.memory\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11674_ _00196_ net467 u_cpu.rf_ram.memory\[44\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07682__A2 _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__A1 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09959__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _04068_ _05172_ _05175_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08631__A1 u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _05130_ _05132_ u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06088__I3 u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10487_ _02862_ _03281_ _05088_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11518__A1 u_cpu.rf_ram.memory\[100\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09187__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12226_ _00740_ net346 u_cpu.rf_ram.memory\[124\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07198__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12157_ _00671_ net79 u_cpu.rf_ram.memory\[131\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10741__A2 _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11108_ u_cpu.rf_ram.memory\[108\]\[1\] _05490_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12088_ _00602_ net72 u_cpu.rf_ram.memory\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout196_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11039_ u_cpu.rf_ram.memory\[106\]\[1\] _05445_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__I u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08698__A1 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06548__I1 u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout363_I net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07370__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06580_ _01915_ _02223_ _01807_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10257__A1 _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout530_I net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08250_ _03500_ _03514_ _03519_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08870__A1 u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07201_ _02769_ _02765_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08181_ _03415_ _03469_ _03474_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09885__I _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07132_ _02709_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10029__C _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08622__A1 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06484__I0 u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07063_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_dbus_dat\[13\] _02665_ _02668_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05918__I _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10980__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06014_ _01610_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07189__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10732__A2 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06400__A3 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07965_ _03326_ _03330_ _03332_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09704_ u_cpu.rf_ram.memory\[115\]\[5\] _04451_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06916_ _02518_ _02531_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _03283_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09125__I _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ u_cpu.rf_ram.memory\[11\]\[5\] _04406_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09350__A2 _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06847_ _01452_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07361__A1 u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06778_ u_cpu.rf_ram.memory\[124\]\[7\] u_cpu.rf_ram.memory\[125\]\[7\] u_cpu.rf_ram.memory\[126\]\[7\]
+ u_cpu.rf_ram.memory\[127\]\[7\] _01706_ _01707_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09566_ _04337_ _04365_ _04368_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08517_ _03053_ _03595_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09497_ u_cpu.rf_ram.memory\[34\]\[1\] _04322_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07113__A1 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10799__A2 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__A1 u_cpu.rf_ram.memory\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _03647_ _03625_ _03648_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08379_ _03596_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ _04816_ _05036_ _05044_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08613__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11390_ u_cpu.rf_ram.memory\[27\]\[2\] _05674_ _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11777__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ u_cpu.cpu.immdec.imm19_12_20\[7\] _04676_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05978__A2 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09169__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _04831_ _04745_ _04932_ _04713_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12011_ _00525_ net56 u_cpu.rf_ram.memory\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout460 net470 net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout471 net473 net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout482 net483 net482 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout493 net494 net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12402__CLK net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10487__A1 _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12913_ _01410_ net196 u_cpu.rf_ram.memory\[100\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12844_ _01341_ net435 u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10239__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07104__A1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12775_ _01272_ net11 u_cpu.rf_ram.memory\[69\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12552__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06394__I _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11726_ _00248_ net210 u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06702__I1 u_cpu.rf_ram.memory\[89\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11657_ _00179_ net403 u_cpu.rf_ram.memory\[46\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _04807_ _05160_ _05165_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08604__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _00110_ net411 u_cpu.rf_ram.memory\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__I0 u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout111_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10539_ _05122_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout209_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A3 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12209_ _00723_ net301 u_cpu.rf_ram.memory\[126\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10714__A2 _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout480_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__A2 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07591__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07750_ u_cpu.rf_ram.memory\[41\]\[0\] _03186_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10312__C _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06701_ _01615_ _02343_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09332__A2 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ _03133_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09420_ u_cpu.rf_ram.memory\[90\]\[3\] _04271_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06632_ u_cpu.rf_ram.memory\[136\]\[5\] u_cpu.rf_ram.memory\[137\]\[5\] u_cpu.rf_ram.memory\[138\]\[5\]
+ u_cpu.rf_ram.memory\[139\]\[5\] _01764_ _01875_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08784__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07894__A2 _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06563_ _02200_ _02202_ _02204_ _02206_ _01717_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09351_ _04171_ _04218_ _04225_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06529__S0 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ _03167_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09282_ _04158_ _04181_ _04184_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout24_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08843__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06494_ _01919_ _02138_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ u_cpu.rf_ram.memory\[66\]\[5\] _03501_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10650__A1 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08164_ u_cpu.rf_ram.memory\[6\]\[4\] _03461_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09399__A2 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10402__A1 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07115_ _02699_ _02696_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _03418_ _03410_ _03419_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08071__A2 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07046_ _02633_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06472__I3 u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06909__A1 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10705__A2 _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12425__CLK net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__A2 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08997_ u_cpu.rf_ram.memory\[134\]\[0\] _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07582__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _03220_ _03314_ _03320_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05983__I2 u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07879_ u_cpu.rf_ram.memory\[4\]\[7\] _03258_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07334__A1 _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12575__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09618_ u_cpu.rf_ram.memory\[8\]\[7\] _04388_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ u_cpu.rf_ram.memory\[101\]\[1\] _05352_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09549_ _04339_ _04353_ _04358_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12560_ _01058_ net308 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08834__A1 u_cpu.rf_ram.memory\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11511_ _03630_ _05742_ _05747_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__I1 _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12491_ _00992_ net237 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11442_ _05310_ _03327_ _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06860__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11197__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _01480_ _02503_ _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10944__A2 _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10324_ _04705_ _04728_ _04962_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07270__B1 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10255_ _04916_ _04917_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09011__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10186_ _04687_ _04854_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07573__A1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11295__I _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout290 net304 net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09314__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06128__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07325__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07876__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__A3 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10180__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11942__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05887__B2 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12827_ _01324_ net107 u_cpu.rf_ram.memory\[86\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout159_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12758_ _01255_ net207 u_cpu.rf_ram.memory\[83\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07628__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08109__I _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07013__I _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10632__A1 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11709_ _00231_ net374 u_cpu.rf_ram.memory\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout326_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12689_ _01186_ net170 u_cpu.rf_ram.memory\[101\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06931__S0 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06852__I u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11188__A2 _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10374__I _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08053__A2 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__I1 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout9 net14 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10935__A2 _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05811__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ _03945_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10699__A1 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ _03628_ _03902_ _03905_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09553__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06367__A2 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12598__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _02927_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08782_ _03861_ _03846_ _03862_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05994_ _01621_ _01627_ _01633_ _01641_ _01642_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07733_ _03139_ _03170_ _03175_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11112__A2 _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07664_ u_cpu.rf_ram.memory\[46\]\[6\] _03122_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05931__I _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09403_ _04260_ _04249_ _04261_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06615_ _01672_ _02258_ _01963_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07595_ _03031_ _03071_ _03080_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06546_ u_cpu.rf_ram.memory\[140\]\[4\] u_cpu.rf_ram.memory\[141\]\[4\] u_cpu.rf_ram.memory\[142\]\[4\]
+ u_cpu.rf_ram.memory\[143\]\[4\] _02101_ _01749_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09334_ u_cpu.rf_ram.memory\[37\]\[7\] _04204_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07619__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08816__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10623__A1 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06477_ u_cpu.rf_ram.memory\[0\]\[4\] u_cpu.rf_ram.memory\[1\]\[4\] u_cpu.rf_ram.memory\[2\]\[4\]
+ u_cpu.rf_ram.memory\[3\]\[4\] _01786_ _01900_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09265_ u_cpu.rf_ram.memory\[124\]\[5\] _04162_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08292__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08216_ _03494_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09196_ _04099_ _04117_ _04125_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11179__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ u_cpu.rf_ram.memory\[75\]\[7\] _03441_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09241__A1 _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08044__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ u_cpu.rf_ram.memory\[77\]\[7\] _03396_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09792__A2 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06150__S1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07029_ _02646_ _02643_ _02639_ _02647_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11815__CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10040_ _04726_ _04630_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09544__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06602__I0 u_cpu.rf_ram.memory\[124\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11965__CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06002__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11991_ _00513_ net420 u_cpu.rf_ram.memory\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11103__A2 _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10942_ u_cpu.rf_ram.memory\[103\]\[6\] _05380_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07858__A2 _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10873_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _05341_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06530__A2 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12612_ _01109_ net444 u_cpu.rf_ram.memory\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08807__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10614__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12543_ _00022_ net252 u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07768__I _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12474_ _00975_ net259 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11425_ u_cpu.rf_ram.memory\[25\]\[0\] _05695_ _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08035__A2 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11356_ _05650_ _02515_ _01461_ _02617_ _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06141__S1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__A1 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ _04728_ _04655_ _04962_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11287_ u_cpu.rf_ram.memory\[111\]\[5\] _05599_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__A2 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13026_ _00088_ net535 u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10238_ _04617_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07546__A1 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11342__A2 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10169_ _04281_ _02627_ _01445_ _02461_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10550__B1 _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout276_I net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout443_I net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12120__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06400_ _01795_ _02033_ _02045_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_91_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _02925_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10605__A1 _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06331_ _01730_ _01977_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10456__I1 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09471__A1 _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08274__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09050_ u_cpu.rf_ram.memory\[132\]\[2\] _04031_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10081__A2 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06262_ u_cpu.rf_ram.memory\[36\]\[2\] u_cpu.rf_ram.memory\[37\]\[2\] u_cpu.rf_ram.memory\[38\]\[2\]
+ u_cpu.rf_ram.memory\[39\]\[2\] _01797_ _01586_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10318__B _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _03326_ _03358_ _03360_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06193_ u_cpu.rf_ram.memory\[112\]\[1\] u_cpu.rf_ram.memory\[113\]\[1\] u_cpu.rf_ram.memory\[114\]\[1\]
+ u_cpu.rf_ram.memory\[115\]\[1\] _01679_ _01840_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09223__A1 _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07085__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _04605_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout91_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11988__CLK net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _03937_ _03927_ _03938_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09526__A2 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__I _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09883_ _02692_ _04526_ _04583_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11333__A2 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ u_cpu.rf_ram.memory\[143\]\[3\] _03893_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08765_ _03844_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05977_ _01483_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _03146_ _03156_ _03163_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _03806_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10844__A1 u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07647_ _03031_ _03107_ _03116_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _03069_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12613__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09317_ _04204_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06529_ u_cpu.rf_ram.memory\[84\]\[4\] u_cpu.rf_ram.memory\[85\]\[4\] u_cpu.rf_ram.memory\[86\]\[4\]
+ u_cpu.rf_ram.memory\[87\]\[4\] _01855_ _02083_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A1 u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08265__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10072__A2 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09248_ u_cpu.rf_ram.memory\[124\]\[1\] _04155_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__S1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08017__A2 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09214__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09179_ _03230_ _03356_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06028__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11210_ _05550_ _05552_ _05554_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07076__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12190_ _00704_ net260 u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10742__I _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ u_cpu.rf_ram.memory\[69\]\[7\] _05500_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05882__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11072_ _05415_ _05458_ _05466_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09517__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11324__A2 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10023_ _04702_ _04704_ _04710_ _04711_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11974_ _00496_ net29 u_cpu.rf_ram.memory\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09043__I _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10835__A1 u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ _05157_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09978__I _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12293__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10856_ _05334_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A2 _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10787_ u_cpu.rf_ram.memory\[95\]\[4\] _05287_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12526_ _01027_ net322 u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06806__A3 _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06362__S1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12457_ _00958_ net252 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09205__A1 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08008__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07067__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _05623_ _05682_ _05685_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12388_ _00889_ net472 u_cpu.rf_ram.memory\[122\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06814__I0 u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11339_ u_cpu.rf_ram.memory\[88\]\[7\] _05619_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06351__B _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09508__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout393_I net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05900_ _01548_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13009_ _00069_ net530 u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06880_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.init_done _02519_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05831_ _01478_ _01455_ _01479_ _01447_ _01481_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11483__I _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08550_ _03673_ _03706_ _03713_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12636__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10320__C _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07501_ _03010_ _03015_ _03017_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10826__A1 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08481_ _03668_ _03663_ _03670_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07432_ _02919_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10827__I _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08247__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07363_ _02903_ u_cpu.rf_ram_if.wdata1_r\[1\] _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11660__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__A1 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09102_ _02907_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06258__A1 _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06314_ _01635_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11251__A1 u_cpu.rf_ram.memory\[110\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09995__A2 _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07294_ _02766_ u_scanchain_local.module_data_in\[68\] _02767_ u_arbiter.i_wb_cpu_dbus_adr\[31\]
+ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06245_ u_cpu.rf_ram.memory\[20\]\[2\] u_cpu.rf_ram.memory\[21\]\[2\] u_cpu.rf_ram.memory\[22\]\[2\]
+ u_cpu.rf_ram.memory\[23\]\[2\] _01891_ _01525_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09033_ _04003_ _04015_ _04021_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11003__A1 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__B1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06176_ _01592_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09747__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07758__A1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11554__A2 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09128__I _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09935_ _03274_ u_arbiter.i_wb_cpu_rdt\[13\] _04626_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06281__I1 u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11306__A2 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12166__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__A2 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09866_ _04572_ _04573_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10365__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08183__A1 _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08817_ u_cpu.rf_ram.memory\[70\]\[5\] _03880_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _04519_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06584__I2 u_cpu.rf_ram.memory\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _03746_ _03832_ _03839_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10817__A1 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08679_ u_cpu.rf_ram.memory\[141\]\[1\] _03796_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08486__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _05232_ _05236_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11490__A1 u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11690_ _00212_ net457 u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10641_ _05183_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10737__I _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11242__A1 _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__B2 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _05137_ _05139_ u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07997__A1 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12311_ _00812_ net487 u_cpu.rf_ram.memory\[35\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07049__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09738__A2 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12242_ _00743_ net358 u_cpu.rf_ram.memory\[123\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11545__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10202__C1 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12509__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12173_ _00687_ net424 u_cpu.rf_ram.memory\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11124_ _05500_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06972__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11055_ _03196_ _05455_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12659__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10006_ _04689_ _04693_ _04695_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A1 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10808__A1 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11957_ _00479_ net23 u_cpu.rf_ram.memory\[54\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11683__CLK net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08477__A2 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06032__S0 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11481__A1 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ u_cpu.rf_ram.memory\[102\]\[0\] _05364_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11888_ _00410_ net270 u_cpu.rf_ram.memory\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout141_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10839_ _05322_ _05312_ _05323_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout239_I net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12039__CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11233__A1 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10036__A2 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__A2 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12509_ _01010_ net188 u_cpu.rf_ram.memory\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout406_I net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06030_ _01583_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06660__A1 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09729__A2 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11536__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_64_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout119 net120 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07981_ u_cpu.rf_ram.memory\[40\]\[4\] _03338_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09720_ u_cpu.rf_ram.memory\[116\]\[3\] _04463_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06932_ _02569_ _02570_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08165__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09901__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ u_cpu.rf_ram.memory\[112\]\[3\] _04418_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06863_ _02498_ _02499_ _02501_ _02502_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_55_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07912__A1 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _03748_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05814_ _01456_ _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09582_ _04376_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06794_ u_cpu.rf_ram.memory\[84\]\[7\] u_cpu.rf_ram.memory\[85\]\[7\] u_cpu.rf_ram.memory\[86\]\[7\]
+ u_cpu.rf_ram.memory\[87\]\[7\] _01684_ _02083_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_83_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06100__I _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08533_ u_cpu.rf_ram.memory\[55\]\[6\] _03698_ _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__A2 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _03577_ _03651_ _03658_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07415_ u_cpu.raddr\[1\] _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08395_ u_cpu.rf_ram.memory\[19\]\[0\] _03610_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10027__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__A2 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07346_ _02876_ u_cpu.rf_ram_if.wen1_r _01438_ u_cpu.rf_ram_if.wen0_r _02895_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06326__S1 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _02630_ _02831_ _02834_ _02835_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08640__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09016_ u_cpu.rf_ram.memory\[134\]\[6\] _04001_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06228_ u_cpu.rf_ram.memory\[128\]\[1\] u_cpu.rf_ram.memory\[129\]\[1\] u_cpu.rf_ram.memory\[130\]\[1\]
+ u_cpu.rf_ram.memory\[131\]\[1\] _01747_ _01875_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06651__B2 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06159_ _01610_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12801__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _02706_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08156__A1 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09849_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _04557_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07903__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12860_ _01357_ net241 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12951__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06010__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11811_ _00333_ net35 u_cpu.rf_ram.memory\[75\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09656__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08459__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12791_ _01288_ net165 u_cpu.rf_ram.memory\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11742_ _00264_ net430 u_cpu.rf_ram.memory\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06945__I _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11673_ _00195_ net466 u_cpu.rf_ram.memory\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06190__I0 u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10624_ u_cpu.rf_ram.memory\[3\]\[1\] _05173_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09959__A2 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10555_ _05109_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08631__A2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06642__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10486_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] _02501_ _03281_
+ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11518__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05996__A3 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12225_ _00739_ net345 u_cpu.rf_ram.memory\[124\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10726__B1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__A1 u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07198__A2 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06245__I1 u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12481__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _00670_ net82 u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11107_ _05468_ _05489_ _05491_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12087_ _00601_ net64 u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11038_ _05399_ _05444_ _05446_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09895__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10151__B _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08698__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06173__A3 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09647__A1 _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12989_ _00047_ net519 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10257__A2 _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout523_I net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07200_ _02724_ _02770_ _02771_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11206__A1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06881__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08180_ u_cpu.rf_ram.memory\[68\]\[2\] _03473_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07131_ _02713_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06804__B _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07062_ _02667_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06013_ u_cpu.rf_ram.memory\[104\]\[0\] u_cpu.rf_ram.memory\[105\]\[0\] u_cpu.rf_ram.memory\[106\]\[0\]
+ u_cpu.rf_ram.memory\[107\]\[0\] _01661_ _01571_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11001__I _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10717__B1 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06936__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10732__A3 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10840__I _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ u_cpu.rf_ram.memory\[40\]\[0\] _03331_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12974__CLK net518 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08138__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05934__I _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09703_ _04438_ _04447_ _04454_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06915_ _02547_ _02548_ _02553_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07895_ u_arbiter.i_wb_cpu_dbus_dat\[3\] u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ u_arbiter.i_wb_cpu_dbus_dat\[1\] _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08689__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09634_ _04075_ _04402_ _04409_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06846_ _02485_ u_cpu.cpu.bne_or_bge _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12204__CLK net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07361__A2 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09565_ u_cpu.rf_ram.memory\[118\]\[1\] _04366_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09638__A1 _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06777_ _02412_ _02414_ _02416_ _02418_ _01577_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_83_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _03679_ _03683_ _03692_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09496_ _04246_ _04321_ _04323_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08447_ u_cpu.rf_ram.memory\[5\]\[7\] _03623_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08861__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06711__I2 u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06872__A1 _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08980__I _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ _03568_ _03597_ _03600_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02514_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08613__A2 _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10340_ _04992_ _04993_ _04941_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _04637_ _04726_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__A1 u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12010_ _00524_ net67 u_cpu.rf_ram.memory\[142\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06005__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout450 net451 net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_94_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout461 net462 net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout472 net476 net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout483 net484 net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout494 net495 net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12912_ _01409_ net196 u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10487__A2 _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12843_ _01340_ net107 u_cpu.rf_ram.memory\[87\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__A1 u_cpu.rf_ram.memory\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10239__A2 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12774_ _01271_ net11 u_cpu.rf_ram.memory\[69\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__A1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07104__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06538__S1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11725_ _00247_ net376 u_cpu.rf_ram.memory\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10197__I _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06863__A1 _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ _00178_ net403 u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11721__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12847__CLK net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10607_ u_cpu.rf_ram.memory\[109\]\[2\] _05164_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10925__I _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ _00109_ net411 u_cpu.rf_ram.memory\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09801__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08604__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06615__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10538_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _05116_ _05118_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12997__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10469_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _05072_
+ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08368__A1 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12208_ _00722_ net301 u_cpu.rf_ram.memory\[126\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10660__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06769__I2 u_cpu.rf_ram.memory\[102\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12139_ _00653_ net77 u_cpu.rf_ram.memory\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07591__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08130__I _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout473_I net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09868__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__B2 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06700_ u_cpu.rf_ram.memory\[92\]\[6\] u_cpu.rf_ram.memory\[93\]\[6\] u_cpu.rf_ram.memory\[94\]\[6\]
+ u_cpu.rf_ram.memory\[95\]\[6\] _02075_ _01619_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07680_ _02920_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08540__A1 u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06631_ _02255_ _02274_ _01475_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ u_cpu.rf_ram.memory\[36\]\[5\] _04221_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06562_ _02006_ _02205_ _01728_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09096__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06529__S1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08301_ _03511_ _03540_ _03549_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ u_cpu.rf_ram.memory\[123\]\[1\] _04182_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06493_ u_cpu.rf_ram.memory\[60\]\[4\] u_cpu.rf_ram.memory\[61\]\[4\] u_cpu.rf_ram.memory\[62\]\[4\]
+ u_cpu.rf_ram.memory\[63\]\[4\] _01617_ _02034_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06854__A1 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08232_ _03346_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10650__A2 _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout17_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _02928_ _03457_ _03463_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05929__I _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07114_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10402__A2 _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ u_cpu.rf_ram.memory\[74\]\[3\] _03416_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07045_ _02657_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13002__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _03994_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07582__A2 _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ u_cpu.rf_ram.memory\[17\]\[3\] _03318_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__B2 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08975__I _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ _02946_ _03260_ _03268_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08531__A1 u_cpu.rf_ram.memory\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _04079_ _04390_ _04398_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06829_ u_arbiter.i_wb_cpu_dbus_we _02468_ u_cpu.cpu.immdec.imm24_20\[0\] _02470_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ u_cpu.rf_ram.memory\[120\]\[2\] _04357_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11744__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09087__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09479_ _04308_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11510_ u_cpu.rf_ram.memory\[100\]\[2\] _05746_ _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12490_ _00991_ net237 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__I1 u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11441_ _05636_ _05695_ _05704_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11894__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06448__I1 u_cpu.rf_ram.memory\[77\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08215__I _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11372_ _05659_ _05661_ _05662_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07259__C _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10323_ _04705_ _04974_ _04975_ _04977_ _04700_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07270__A1 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10254_ u_cpu.cpu.immdec.imm30_25\[4\] _04880_ _04905_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _04913_ _04683_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__10157__A1 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09011__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__S0 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10185_ _04743_ _04713_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08770__A1 _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout280 net284 net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout291 net293 net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06208__S0 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08885__I _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10180__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05887__A2 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12826_ _01323_ net118 u_cpu.rf_ram.memory\[86\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09078__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12757_ _01254_ net186 u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11708_ _00230_ net388 u_cpu.rf_ram.memory\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10632__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12688_ _01185_ net194 u_cpu.rf_ram.memory\[101\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11639_ _00161_ net163 u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13025__CLK net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout319_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05811__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11617__CLK net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ u_cpu.rf_ram.memory\[14\]\[1\] _03903_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07185__B _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10323__C _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07801_ _03217_ _03212_ _03219_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ u_cpu.rf_ram.memory\[73\]\[7\] _03844_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05993_ _01488_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07732_ u_cpu.rf_ram.memory\[51\]\[2\] _03174_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11767__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07663_ _03027_ _03119_ _03126_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10320__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ u_cpu.rf_ram.memory\[91\]\[5\] _04254_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06614_ u_cpu.rf_ram.memory\[88\]\[5\] u_cpu.rf_ram.memory\[89\]\[5\] u_cpu.rf_ram.memory\[90\]\[5\]
+ u_cpu.rf_ram.memory\[91\]\[5\] _01961_ _01674_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07594_ u_cpu.rf_ram.memory\[80\]\[7\] _03069_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09333_ _04174_ _04206_ _04214_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06545_ _02188_ _02189_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08816__A2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10623__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _04170_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06476_ _02011_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _03494_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09195_ u_cpu.rf_ram.memory\[127\]\[6\] _04120_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ _03424_ _03443_ _03451_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10387__A1 u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09241__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ _03350_ _03398_ _03406_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07028_ _02492_ _02612_ _02635_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05802__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10514__B _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06438__S0 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12542__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08979_ _03930_ _03982_ _03985_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11990_ _00512_ net420 u_cpu.rf_ram.memory\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07307__A2 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10941_ _05324_ _05377_ _05384_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10311__A1 _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10872_ _05343_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07114__I u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12611_ _01108_ net444 u_cpu.rf_ram.memory\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08807__A2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12542_ _01043_ net318 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06818__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09480__A2 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12473_ _00974_ net237 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11424_ _05693_ _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12072__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10378__A1 u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__A2 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11355_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07794__A2 _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _04747_ _04662_ _04630_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08991__A1 u_cpu.rf_ram.memory\[135\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11286_ _05562_ _05595_ _05602_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13025_ _00087_ net535 u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10237_ _04898_ _04900_ _04824_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10168_ _01457_ _04677_ _04840_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10550__B2 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10099_ _04691_ _04706_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_43_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout171_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout269_I net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12809_ _01306_ net111 u_cpu.rf_ram.memory\[85\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout436_I net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ u_cpu.rf_ram.memory\[72\]\[2\] u_cpu.rf_ram.memory\[73\]\[2\] u_cpu.rf_ram.memory\[74\]\[2\]
+ u_cpu.rf_ram.memory\[75\]\[2\] _01867_ _01732_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10605__A2 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12415__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06261_ _01899_ _01903_ _01905_ _01907_ _01578_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07482__A1 _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__A2 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08000_ u_cpu.rf_ram.memory\[119\]\[0\] _03359_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__C _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06192_ _01585_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09223__A2 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07234__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11030__A2 _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12565__CLK net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07085__I1 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07785__A2 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08982__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ _04629_ _04642_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06531__C _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08902_ u_cpu.rf_ram.memory\[39\]\[4\] _03933_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09882_ u_arbiter.i_wb_cpu_rdt\[31\] _04492_ _04574_ _02478_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout84_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A1 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07537__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06103__I _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _03850_ _03889_ _03894_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _03738_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05976_ u_cpu.rf_ram.memory\[56\]\[0\] u_cpu.rf_ram.memory\[57\]\[0\] u_cpu.rf_ram.memory\[58\]\[0\]
+ u_cpu.rf_ram.memory\[59\]\[0\] _01623_ _01624_ _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05942__I u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ u_cpu.rf_ram.memory\[44\]\[5\] _03159_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08695_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07646_ u_cpu.rf_ram.memory\[42\]\[7\] _03105_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10844__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07170__B1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ _03069_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09316_ _02960_ _03104_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06528_ _01852_ _02172_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07473__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _04157_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06459_ _01758_ _02104_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12908__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09178_ _04101_ _04105_ _04114_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06028__A2 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08129_ _03440_ _03197_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08973__A1 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _05484_ _05502_ _05510_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11932__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10780__A1 u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__C _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11071_ u_cpu.rf_ram.memory\[107\]\[6\] _05461_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05882__S1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10022_ _04693_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__I u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11973_ _00495_ net29 u_cpu.rf_ram.memory\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06339__I0 u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10924_ _05328_ _05364_ _05373_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10835__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06503__A3 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10855_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _05331_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10786_ _05209_ _05283_ _05289_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10599__A1 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__A1 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12525_ _01026_ net322 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09994__I _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12456_ _00957_ net253 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09205__A2 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11407_ u_cpu.rf_ram.memory\[26\]\[1\] _05683_ _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07216__A1 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10933__I _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__A2 _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12387_ _00888_ net473 u_cpu.rf_ram.memory\[122\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08964__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11338_ _02950_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10771__A1 u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11269_ u_cpu.rf_ram.memory\[86\]\[6\] _05587_ _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13008_ _00068_ net530 u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout386_I net409 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05830_ _01440_ _01480_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07500_ u_cpu.rf_ram.memory\[20\]\[0\] _03016_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ u_cpu.rf_ram.memory\[57\]\[2\] _03669_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07298__A4 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07431_ _02969_ _02966_ _02970_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11805__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06807__B _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07362_ _02901_ _02908_ _02910_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09101_ _04011_ _04052_ _04061_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06313_ _01693_ _01959_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11251__A2 _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07293_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _02844_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09995__A3 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09032_ u_cpu.rf_ram.memory\[133\]\[3\] _04019_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06244_ _01720_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11955__CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07207__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10843__I _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11003__A2 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06175_ _01646_ _01822_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05937__I _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06261__C _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _02705_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08707__A1 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ u_arbiter.i_wb_cpu_rdt\[24\] _04495_ _04521_ u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10514__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10365__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09380__A1 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08183__A2 _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08816_ _03855_ _03876_ _03883_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06194__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ u_arbiter.i_wb_cpu_rdt\[5\] _04512_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09144__I _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ u_cpu.rf_ram.memory\[72\]\[4\] _03836_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06584__I3 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05959_ _01607_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__A1 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10278__B1 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10817__A2 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08678_ _03730_ _03795_ _03797_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07694__A1 u_cpu.rf_ram.memory\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07629_ _03105_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11490__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12730__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10640_ _05183_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07446__A1 u_cpu.rf_ram.memory\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__A2 _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11242__A2 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _05141_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12310_ _00811_ net467 u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07997__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11996__D _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__A1 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12241_ _00742_ net361 u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07049__I1 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05847__I _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12172_ _00686_ net425 u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08223__I _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10202__C2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12110__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11123_ _02960_ _03395_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11054_ _05157_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10505__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10702__B _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10005_ _03277_ _04694_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12260__CLK net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A1 u_cpu.rf_ram.memory\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11828__CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10808__A2 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11956_ _00478_ net23 u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10928__I _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10907_ _05362_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06032__S1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11481__A2 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11887_ _00409_ net89 u_cpu.rf_ram.memory\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10838_ u_cpu.rf_ram.memory\[28\]\[4\] _05318_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11978__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A1 u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11233__A2 _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10769_ u_cpu.rf_ram.memory\[94\]\[5\] _05275_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout134_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10864__S _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12508_ _01009_ net172 u_cpu.rf_ram.memory\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10992__A1 u_cpu.rf_ram.memory\[99\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10663__I _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12439_ _00940_ net246 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout301_I net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08937__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__A1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07980_ _03343_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_68_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12603__CLK net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.bufreg.lsb\[1\]
+ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08165__A2 _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09650_ _04339_ _04414_ _04419_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06862_ u_cpu.cpu.decode.op26 _01447_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08601_ _02937_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05813_ _01458_ _01459_ _01438_ _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_94_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09581_ _04376_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06793_ _01678_ _02434_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__A1 u_cpu.rf_ram.memory\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08532_ _03675_ _03695_ _03702_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout47_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07676__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ u_cpu.rf_ram.memory\[58\]\[5\] _03654_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11472__A2 _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07414_ _02885_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.raddr\[0\] u_cpu.rf_ram_if.rcnt\[2\]
+ _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ _03608_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07428__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ u_cpu.cpu.immdec.imm11_7\[4\] _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _02757_ _02766_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09015_ _03751_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12133__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06227_ _01748_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08928__A1 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06158_ u_cpu.rf_ram.memory\[44\]\[1\] u_cpu.rf_ram.memory\[45\]\[1\] u_cpu.rf_ram.memory\[46\]\[1\]
+ u_cpu.rf_ram.memory\[47\]\[1\] _01805_ _01608_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10735__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06089_ _01484_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07882__I _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12283__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09917_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _04604_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08156__A2 _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09353__A1 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09848_ _04558_ _04561_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11160__A1 u_cpu.rf_ram.memory\[84\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07903__A2 _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06262__S1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _04505_ _04507_ _04491_ _04508_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11810_ _00332_ net126 u_cpu.rf_ram.memory\[76\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12790_ _01287_ net73 u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09602__I _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _00263_ net435 u_cpu.rf_ram.memory\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07667__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11672_ _00194_ net466 u_cpu.rf_ram.memory\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07122__I _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10623_ _04062_ _05172_ _05174_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06890__A2 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10554_ _05131_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08092__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10974__A1 _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06642__A2 _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10485_ _05087_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09049__I _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08919__A1 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12224_ _00738_ net350 u_cpu.rf_ram.memory\[124\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12626__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10726__A1 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10726__B2 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12155_ _00669_ net80 u_cpu.rf_ram.memory\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__I2 u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__I _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ u_cpu.rf_ram.memory\[108\]\[0\] _05490_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12086_ _00600_ net64 u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11650__CLK net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09344__A1 u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08147__A2 _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ u_cpu.rf_ram.memory\[106\]\[0\] _05445_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12776__CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09895__A2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12006__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09647__A2 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12988_ _00046_ net517 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09512__I _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout251_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11454__A2 _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11939_ _00461_ net68 u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout349_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08128__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11206__A2 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12156__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout516_I net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06881__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07967__I _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07130_ _02695_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11489__I _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10965__A1 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ u_arbiter.i_wb_cpu_rdt\[15\] u_arbiter.i_wb_cpu_dbus_dat\[12\] _02665_ _02667_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07830__A1 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06633__A2 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10017__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06012_ _01605_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__A1 _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08386__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ _03329_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09335__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08138__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09702_ u_cpu.rf_ram.memory\[115\]\[4\] _04451_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06914_ _02549_ _02533_ _02551_ _02552_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07894_ _03280_ _03281_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11142__A1 _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09633_ u_cpu.rf_ram.memory\[11\]\[4\] _04406_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07897__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06845_ _01451_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06111__I _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09564_ _04332_ _04365_ _04367_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06776_ _02055_ _02417_ _02058_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09638__A2 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05950__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ u_cpu.rf_ram.memory\[56\]\[7\] _03681_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11445__A2 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ u_cpu.rf_ram.memory\[34\]\[0\] _04322_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _03646_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__A2 _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08377_ u_cpu.rf_ram.memory\[60\]\[1\] _03598_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10256__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07328_ _02514_ _01458_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12649__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08074__A1 u_cpu.rf_ram.memory\[77\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _02757_ _02818_ _02820_ _02766_ _02821_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06624__A2 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06475__I2 u_cpu.rf_ram.memory\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06180__S0 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10270_ _04700_ _04930_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10708__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__A2 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06730__B _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11381__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout440 net449 net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout451 net510 net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout462 net463 net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout473 net476 net473 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__12029__CLK net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout484 net494 net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout495 net509 net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12911_ _01408_ net175 u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07888__A1 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12842_ _01339_ net118 u_cpu.rf_ram.memory\[87\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06560__A1 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09629__A2 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07053__S _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11436__A2 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12179__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10239__A3 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12773_ _01270_ net12 u_cpu.rf_ram.memory\[69\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__A2 _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11724_ _00246_ net375 u_cpu.rf_ram.memory\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11655_ _00177_ net405 u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net81 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06905__B u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 net92 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_10606_ _05159_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08065__A1 u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11586_ _00108_ net411 u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09801__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _05121_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07812__A1 u_cpu.rf_ram.memory\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _05076_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08368__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12207_ _00721_ net299 u_cpu.rf_ram.memory\[126\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10399_ _04805_ _05035_ _05038_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _00652_ net82 u_cpu.rf_ram.memory\[134\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout299_I net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12069_ _00583_ net58 u_cpu.rf_ram.memory\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09868__A2 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout466_I net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06630_ _01958_ _02264_ _02273_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08540__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09242__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06561_ u_cpu.rf_ram.memory\[16\]\[5\] u_cpu.rf_ram.memory\[17\]\[5\] u_cpu.rf_ram.memory\[18\]\[5\]
+ u_cpu.rf_ram.memory\[19\]\[5\] _02007_ _01518_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11427__A2 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ u_cpu.rf_ram.memory\[29\]\[7\] _03538_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _04152_ _04181_ _04183_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06492_ _02130_ _02132_ _02134_ _02136_ _01665_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08231_ _03505_ _03495_ _03506_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06854__A2 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__B _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08162_ u_cpu.rf_ram.memory\[6\]\[3\] _03461_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08056__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07113_ _02630_ u_scanchain_local.module_data_in\[38\] _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11696__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ _03340_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06162__S0 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ u_arbiter.i_wb_cpu_rdt\[8\] u_arbiter.i_wb_cpu_dbus_dat\[5\] _02652_ _02657_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09556__A1 u_cpu.rf_ram.memory\[120\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08359__A2 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10166__A2 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08995_ _03994_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ _03217_ _03314_ _03319_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ u_cpu.rf_ram.memory\[4\]\[6\] _03263_ _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12321__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ u_cpu.rf_ram.memory\[8\]\[6\] _04393_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06828_ u_arbiter.i_wb_cpu_dbus_we _02467_ _02468_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_55_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11418__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _04352_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06759_ _01667_ _02400_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08295__A1 _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ _04251_ _04309_ _04312_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12471__CLK net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ _02926_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11440_ u_cpu.rf_ram.memory\[25\]\[7\] _05693_ _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08047__A1 u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10247__B _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11371_ _02511_ _05661_ _04234_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06448__I2 u_cpu.rf_ram.memory\[78\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _04958_ _04822_ _04889_ _04976_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_50_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06016__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10253_ _04861_ _04912_ _04915_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05855__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _04729_ _04795_ _04851_ _04852_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06456__S1 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout270 net272 net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout281 net283 net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout292 net293 net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06208__S1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A2 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05804__B _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12825_ _01322_ net111 u_cpu.rf_ram.memory\[86\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12756_ _01253_ net186 u_cpu.rf_ram.memory\[83\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11707_ _00229_ net388 u_cpu.rf_ram.memory\[48\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06687__I2 u_cpu.rf_ram.memory\[106\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06836__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12687_ _01184_ net194 u_cpu.rf_ram.memory\[101\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06635__B _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08038__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11638_ _00160_ net163 u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09786__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11569_ _04234_ u_cpu.rf_ram_if.rreq_r _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09538__A1 u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10671__I _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05811__A3 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08210__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10699__A3 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12344__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07800_ u_cpu.rf_ram.memory\[48\]\[2\] _03218_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08780_ _03754_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05992_ _01634_ _01639_ _01640_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06772__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__I _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07731_ _03169_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09710__A1 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A2 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07662_ u_cpu.rf_ram.memory\[46\]\[5\] _03122_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06524__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12494__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06613_ _01615_ _02256_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09401_ _04170_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _03029_ _03071_ _03079_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06544_ u_cpu.rf_ram.memory\[136\]\[4\] u_cpu.rf_ram.memory\[137\]\[4\] u_cpu.rf_ram.memory\[138\]\[4\]
+ u_cpu.rf_ram.memory\[139\]\[4\] _01747_ _01875_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09332_ u_cpu.rf_ram.memory\[37\]\[6\] _04209_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__A1 _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09263_ _02937_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06475_ u_cpu.rf_ram.memory\[4\]\[4\] u_cpu.rf_ram.memory\[5\]\[4\] u_cpu.rf_ram.memory\[6\]\[4\]
+ u_cpu.rf_ram.memory\[7\]\[4\] _01782_ _01897_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10846__I _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08214_ _02891_ _03087_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08029__A1 u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09194_ _04097_ _04117_ _04124_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07220__I _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10067__B _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ u_cpu.rf_ram.memory\[75\]\[6\] _03446_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08076_ u_cpu.rf_ram.memory\[77\]\[6\] _03401_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ u_arbiter.i_wb_cpu_rdt\[2\] _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_122_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11336__A1 u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09147__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06438__S1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08752__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08978_ u_cpu.rf_ram.memory\[135\]\[1\] _03983_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11711__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07929_ u_cpu.rf_ram.memory\[16\]\[4\] _03306_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09701__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10940_ u_cpu.rf_ram.memory\[103\]\[5\] _05380_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__I1 u_cpu.rf_ram.memory\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _05341_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11861__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12987__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12610_ _01107_ net443 u_cpu.rf_ram.memory\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10075__A1 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11999__D _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__I _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06818__A2 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12541_ _01042_ net318 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08226__I _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12217__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12472_ _00973_ net279 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09768__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _05693_ _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11354_ _05642_ _05641_ _05649_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08440__A1 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12367__CLK net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10305_ _04902_ _04727_ _04932_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08991__A2 _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12623__D _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11285_ u_cpu.rf_ram.memory\[111\]\[4\] _05599_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11327__A1 u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10236_ _04828_ _04899_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13024_ _00086_ net535 u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08743__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _04759_ _04820_ _04837_ _04839_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06754__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10550__A2 _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10098_ _04709_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout164_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12808_ _01305_ net112 u_cpu.rf_ram.memory\[85\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10066__A1 _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10666__I _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout331_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12739_ _01236_ net121 u_cpu.rf_ram.memory\[105\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout429_I net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06260_ _01567_ _01906_ _01792_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06285__A3 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08136__I _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _01836_ _01838_ _01676_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__S0 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07975__I _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08431__A1 u_cpu.rf_ram.memory\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09950_ _04627_ _04631_ _04641_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_89_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11318__A1 _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11734__CLK net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _03745_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09881_ _02690_ _04526_ _04524_ _02692_ _04582_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08832_ u_cpu.rf_ram.memory\[143\]\[2\] _03893_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10541__A2 _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08763_ _03848_ _03845_ _03849_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05975_ _01592_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10350__B _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07714_ _03144_ _03155_ _03162_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08694_ _03152_ _03370_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ _03029_ _03107_ _03115_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07170__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ _02899_ _03068_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10057__A1 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06527_ u_cpu.rf_ram.memory\[80\]\[4\] u_cpu.rf_ram.memory\[81\]\[4\] u_cpu.rf_ram.memory\[82\]\[4\]
+ u_cpu.rf_ram.memory\[83\]\[4\] _01584_ _01965_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09998__A1 _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09315_ _04177_ _04194_ _04203_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10576__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05859__I0 u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06458_ u_cpu.rf_ram.memory\[136\]\[3\] u_cpu.rf_ram.memory\[137\]\[3\] u_cpu.rf_ram.memory\[138\]\[3\]
+ u_cpu.rf_ram.memory\[139\]\[3\] _01759_ _01760_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09246_ _02912_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07473__A2 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08670__A1 u_cpu.rf_ram.memory\[142\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09177_ u_cpu.rf_ram.memory\[128\]\[7\] _04103_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06389_ u_cpu.rf_ram.memory\[60\]\[3\] u_cpu.rf_ram.memory\[61\]\[3\] u_cpu.rf_ram.memory\[62\]\[3\]
+ u_cpu.rf_ram.memory\[63\]\[3\] _01617_ _02034_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11557__A1 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08128_ _03086_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07225__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ _03086_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10017__S _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__A2 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11070_ _05413_ _05458_ _05465_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10021_ _04638_ _04705_ _04706_ _04709_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_27_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08725__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09922__A1 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10532__A2 _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11356__B _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10260__B _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13015__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11972_ _00494_ net28 u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10923_ u_cpu.rf_ram.memory\[102\]\[7\] _05362_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__S0 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10854_ _05333_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07061__S _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10048__A1 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11607__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10785_ u_cpu.rf_ram.memory\[95\]\[3\] _05287_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06347__S0 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10599__A2 _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12524_ _01025_ net322 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12455_ _00956_ net252 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07795__I _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11548__A1 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11406_ _05618_ _05682_ _05684_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11757__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12386_ _00887_ net471 u_cpu.rf_ram.memory\[122\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__A1 _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11337_ _05634_ _05621_ _05635_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06814__I2 u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06975__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10771__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11268_ _05564_ _05584_ _05591_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13007_ _00067_ net528 u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10219_ u_cpu.cpu.immdec.imm30_25\[1\] _04882_ _04884_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11199_ u_cpu.rf_ram.memory\[10\]\[5\] _05543_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout281_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout379_I net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__I _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ u_cpu.rf_ram.memory\[21\]\[1\] _02967_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__I _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ u_cpu.rf_ram.memory\[82\]\[0\] _02909_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12532__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06312_ u_cpu.rf_ram.memory\[92\]\[2\] u_cpu.rf_ram.memory\[93\]\[2\] u_cpu.rf_ram.memory\[94\]\[2\]
+ u_cpu.rf_ram.memory\[95\]\[2\] _01694_ _01847_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09100_ u_cpu.rf_ram.memory\[130\]\[7\] _04050_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08652__A1 u_cpu.rf_ram.memory\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07292_ _02842_ _02847_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09031_ _04000_ _04015_ _04020_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06243_ _01467_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11539__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06174_ u_cpu.rf_ram.memory\[100\]\[1\] u_cpu.rf_ram.memory\[101\]\[1\] u_cpu.rf_ram.memory\[102\]\[1\]
+ u_cpu.rf_ram.memory\[103\]\[1\] _01647_ _01648_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08404__A1 u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12682__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10345__B _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10211__A1 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09933_ _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06114__I _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06281__I3 u_cpu.rf_ram.memory\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08707__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09864_ u_arbiter.i_wb_cpu_dbus_dat\[25\] _04524_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06718__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10514__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ u_cpu.rf_ram.memory\[70\]\[4\] _03880_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _04520_ _04522_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__A1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06194__A2 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08746_ _03743_ _03832_ _03838_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05958_ _01591_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10278__A1 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10278__B2 _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05889_ _01537_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10817__A3 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08677_ u_cpu.rf_ram.memory\[141\]\[0\] _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06577__S0 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _03102_ _03104_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07694__A2 _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07559_ u_cpu.rf_ram.memory\[7\]\[1\] _03057_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10570_ _02800_ _05137_ _05139_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08643__A1 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09229_ u_cpu.rf_ram.memory\[125\]\[3\] _04144_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12240_ _00741_ net361 u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06257__I0 u_cpu.rf_ram.memory\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12171_ _00685_ net424 u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10202__B2 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06957__A1 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10753__A2 _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _05486_ _05490_ _05499_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ _05417_ _05445_ _05454_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05863__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10505__A2 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12405__CLK net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10004_ _04612_ _04618_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A2 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10269__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _00477_ net23 u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06568__S0 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12555__CLK net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _05362_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__S _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07685__A2 _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11886_ _00408_ net89 u_cpu.rf_ram.memory\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10837_ _05211_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10768_ _05212_ _05271_ _05278_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12507_ _01008_ net176 u_cpu.rf_ram.memory\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout127_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ _04891_ _04654_ _04665_ _04762_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06740__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10992__A2 _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12438_ _00939_ net246 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12369_ _00870_ net422 u_cpu.rf_ram.memory\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10744__A2 _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout496_I net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06930_ _02491_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\] _02486_ _02569_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12085__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06861_ _02500_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08600_ _03746_ _03732_ _03747_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05812_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06792_ u_cpu.rf_ram.memory\[80\]\[7\] u_cpu.rf_ram.memory\[81\]\[7\] u_cpu.rf_ram.memory\[82\]\[7\]
+ u_cpu.rf_ram.memory\[83\]\[7\] _01584_ _01586_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_83_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09580_ _03182_ _04179_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__A2 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08531_ u_cpu.rf_ram.memory\[55\]\[5\] _03698_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06559__S0 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08462_ _03575_ _03650_ _03657_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07676__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__A1 u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11922__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _02906_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08393_ _03608_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11015__I _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ u_cpu.cpu.immdec.imm11_7\[2\] _02892_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08625__A1 u_cpu.rf_ram.memory\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07428__A2 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06109__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07275_ _02832_ _02827_ _02833_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06731__S0 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10983__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06226_ _01846_ _01873_ _01743_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09014_ _04007_ _03996_ _04008_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06239__I0 u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ _01605_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10735__A2 _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06088_ u_cpu.rf_ram.memory\[76\]\[0\] u_cpu.rf_ram.memory\[77\]\[0\] u_cpu.rf_ram.memory\[78\]\[0\]
+ u_cpu.rf_ram.memory\[79\]\[0\] _01515_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _04607_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09847_ u_arbiter.i_wb_cpu_rdt\[18\] _04559_ _04560_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07364__A1 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12578__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09778_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _04501_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08729_ u_cpu.rf_ram.memory\[13\]\[5\] _03824_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _00262_ net433 u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A1 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07403__I _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11671_ _00193_ net466 u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__I2 u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10622_ u_cpu.rf_ram.memory\[3\]\[0\] _05173_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08616__A1 u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06019__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10553_ _02769_ _05130_ _05125_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08092__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05858__I _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06722__S0 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10484_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _05086_ _05078_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06493__I3 u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08919__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12223_ _00737_ net344 u_cpu.rf_ram.memory\[124\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09041__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__B1 _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__A2 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12154_ _00668_ net82 u_cpu.rf_ram.memory\[132\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09592__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06245__I3 u_cpu.rf_ram.memory\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11105_ _05488_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12085_ _00599_ net63 u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09344__A2 _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11036_ _05443_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06402__I0 u_cpu.rf_ram.memory\[100\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11945__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12987_ _00045_ net516 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08855__A1 u_cpu.rf_ram.memory\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11938_ _00460_ net37 u_cpu.rf_ram.memory\[57\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout244_I net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11869_ _00391_ net166 u_cpu.rf_ram.memory\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout411_I net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10414__A1 _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout509_I net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09280__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__S0 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ _02666_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07830__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06484__I3 u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ _01659_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06092__C _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07983__I _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10717__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11390__A2 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ _03329_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09701_ _04436_ _04447_ _04453_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06913_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02544_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07893_ _02519_ _02525_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07346__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11142__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09632_ _04073_ _04402_ _04408_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06844_ _01463_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12870__CLK net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__I _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09563_ u_cpu.rf_ram.memory\[118\]\[0\] _04366_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06775_ u_cpu.rf_ram.memory\[104\]\[7\] u_cpu.rf_ram.memory\[105\]\[7\] u_cpu.rf_ram.memory\[106\]\[7\]
+ u_cpu.rf_ram.memory\[107\]\[7\] _02056_ _01624_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08514_ _03677_ _03683_ _03691_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09494_ _04320_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _02950_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12100__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08376_ _03563_ _03597_ _03599_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07327_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08074__A2 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06704__S0 _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07258_ _02819_ _02812_ _02783_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06180__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06209_ _01711_ _01856_ _01715_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11818__CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07189_ _02634_ _02761_ _02762_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout430 net434 net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout441 net443 net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09326__A2 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11968__CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout452 net460 net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout463 net469 net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout474 net475 net474 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07337__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout485 net489 net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout496 net498 net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_12910_ _01407_ net175 u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07888__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12841_ _01338_ net114 u_cpu.rf_ram.memory\[87\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08229__I _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08837__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12772_ _01269_ net12 u_cpu.rf_ram.memory\[69\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _00245_ net375 u_cpu.rf_ram.memory\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11654_ _00176_ net401 u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout70 net75 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout81 net83 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10605_ _04805_ _05160_ _05163_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08065__A2 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11585_ _00107_ net411 u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10536_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _05116_ _05118_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09014__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _05072_
+ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _00720_ net298 u_cpu.rf_ram.memory\[126\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09565__A2 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07576__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ u_cpu.rf_ram.memory\[31\]\[1\] _05036_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06640__C _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12137_ _00651_ net62 u_cpu.rf_ram.memory\[134\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10580__B1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12068_ _00582_ net59 u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout194_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07328__A1 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11019_ u_cpu.rf_ram.memory\[105\]\[1\] _05433_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout361_I net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06551__A2 _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout459_I net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _01890_ _02203_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08828__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ _01915_ _02135_ _01807_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08230_ u_cpu.rf_ram.memory\[66\]\[4\] _03501_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12273__CLK net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _02921_ _03457_ _03462_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09253__A1 u_cpu.rf_ram.memory\[124\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08056__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10938__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06067__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__A1 u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07112_ _02694_ _02697_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08092_ _03415_ _03410_ _03417_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06162__S1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07043_ _02656_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09005__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09556__A2 _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__I _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07567__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06614__I0 u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ _03369_ _03454_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07945_ u_cpu.rf_ram.memory\[17\]\[2\] _03318_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07319__A1 _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11115__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ _02940_ _03260_ _03267_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05961__I _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ _04077_ _04390_ _04397_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10579__I _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06827_ u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.decode.opcode\[0\] u_cpu.cpu.decode.opcode\[1\]
+ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05976__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _04337_ _04353_ _04356_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08819__A1 u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06758_ u_cpu.rf_ram.memory\[60\]\[7\] u_cpu.rf_ram.memory\[61\]\[7\] u_cpu.rf_ram.memory\[62\]\[7\]
+ u_cpu.rf_ram.memory\[63\]\[7\] _01668_ _02034_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12616__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ u_cpu.rf_ram.memory\[35\]\[1\] _04310_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08295__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09492__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06689_ _02325_ _02327_ _02329_ _02331_ _01577_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_52_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08428_ _03631_ _03624_ _03633_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__I3 u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11640__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__A2 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09244__A1 u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08359_ u_cpu.rf_ram.memory\[61\]\[2\] _03588_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12766__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10929__A2 _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11051__A1 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11370_ _02502_ _04232_ _05660_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06448__I3 u_cpu.rf_ram.memory\[79\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _04645_ _04745_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11790__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10252_ _04687_ _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11359__B _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07558__A1 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10183_ _04794_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10562__B1 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12146__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout260 net262 net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11106__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__A2 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout271 net272 net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout282 net283 net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__B1 _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout293 net297 net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__05871__I _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__I _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__C _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__A1 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06533__A2 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12824_ _01321_ net113 u_cpu.rf_ram.memory\[86\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12296__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10617__A1 u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12755_ _01252_ net116 u_cpu.rf_ram.memory\[107\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07798__I _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11290__A1 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11706_ _00228_ net296 u_cpu.rf_ram.memory\[48\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12686_ _01183_ net194 u_cpu.rf_ram.memory\[101\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06687__I3 u_cpu.rf_ram.memory\[107\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11637_ _00159_ net190 u_cpu.rf_ram.memory\[80\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08038__A2 _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11042__A1 u_cpu.rf_ram.memory\[106\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06207__I _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11568_ _05780_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07797__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ _05110_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout207_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11499_ _03643_ _05731_ _05739_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08210__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10553__B1 _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10699__A4 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ _01595_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06772__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07730_ _03137_ _03170_ _03173_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12639__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07661_ _03025_ _03118_ _03125_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09710__A2 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06524__A2 _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09400_ _04258_ _04248_ _04259_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06612_ u_cpu.rf_ram.memory\[92\]\[5\] u_cpu.rf_ram.memory\[93\]\[5\] u_cpu.rf_ram.memory\[94\]\[5\]
+ u_cpu.rf_ram.memory\[95\]\[5\] _02075_ _01847_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ u_cpu.rf_ram.memory\[80\]\[6\] _03074_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__A1 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09331_ _04171_ _04206_ _04213_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06543_ _01538_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08277__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12789__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11281__A1 u_cpu.rf_ram.memory\[111\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout22_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09262_ _04168_ _04154_ _04169_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06474_ _02112_ _02114_ _02116_ _02118_ _01717_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08213_ _03325_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08029__A2 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ u_cpu.rf_ram.memory\[127\]\[5\] _04120_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11033__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ _03422_ _03443_ _03450_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06135__S1 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07788__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08075_ _03347_ _03398_ _03405_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05956__I _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07026_ _02642_ _02643_ _02645_ _02639_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09529__A2 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__I _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12169__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__A2 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10544__B1 _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08201__A2 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ _03925_ _03982_ _03984_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06763__A2 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07928_ _03220_ _03302_ _03308_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10147__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10847__A1 u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09701__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ _03036_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06366__I2 u_cpu.rf_ram.memory\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07712__A1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10870_ _05342_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ u_cpu.rf_ram.memory\[117\]\[4\] _04340_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09465__A1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11272__A1 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12540_ _01041_ net318 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05877__I1 u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12471_ _00972_ net475 u_cpu.rf_ram.memory\[114\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11422_ _05310_ _03183_ _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06027__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09768__A2 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11353_ _05641_ _05648_ _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05866__I _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07059__S _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09338__I _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06451__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _04931_ _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08242__I _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11284_ _05560_ _05595_ _05601_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11327__A2 _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13023_ _00085_ net535 u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10235_ _04679_ _04641_ _04829_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06203__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ _04776_ _04838_ _04695_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10721__B _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _04650_ _04779_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10838__A1 u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11686__CLK net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12931__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10012__I _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12807_ _01304_ net119 u_cpu.rf_ram.memory\[85\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10947__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout157_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09456__A1 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08259__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10999_ u_cpu.rf_ram.memory\[79\]\[1\] _05421_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06646__B _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__A2 _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12738_ _01235_ net121 u_cpu.rf_ram.memory\[105\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10168__B _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10883__S _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09208__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12669_ _01166_ net47 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout324_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06190_ u_cpu.rf_ram.memory\[120\]\[1\] u_cpu.rf_ram.memory\[121\]\[1\] u_cpu.rf_ram.memory\[122\]\[1\]
+ u_cpu.rf_ram.memory\[123\]\[1\] _01673_ _01837_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__S1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12311__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08900_ _03935_ _03927_ _03936_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09880_ u_arbiter.i_wb_cpu_rdt\[30\] _04491_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10526__B1 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07991__I _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12461__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08831_ _03888_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ u_cpu.rf_ram.memory\[73\]\[1\] _03846_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05974_ _01548_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07713_ u_cpu.rf_ram.memory\[44\]\[4\] _03159_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10829__A1 _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08693_ _03755_ _03796_ _03805_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07644_ u_cpu.rf_ram.memory\[42\]\[6\] _03110_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10857__I _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07575_ _03067_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09447__A1 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ u_cpu.rf_ram.memory\[38\]\[7\] _04192_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06526_ _01672_ _02170_ _01963_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10057__A2 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09998__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05859__I1 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09245_ _04152_ _04154_ _04156_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06457_ _01752_ _02102_ _01485_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08670__A2 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09176_ _04099_ _04105_ _04113_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06388_ _01618_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11557__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__I0 u_cpu.rf_ram.memory\[128\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08127_ _03426_ _03430_ _03439_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06433__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ _03353_ _03385_ _03394_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12804__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07009_ _02627_ _02625_ _02631_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10020_ _04708_ _04691_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07933__A1 u_cpu.rf_ram.memory\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06292__S0 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11356__C _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11971_ _00493_ net28 u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09686__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08489__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06339__I2 u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11493__A1 _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10922_ _05326_ _05364_ _05372_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__S1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _05331_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11245__A1 u_cpu.rf_ram.memory\[110\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09989__A2 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10784_ _05205_ _05283_ _05288_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06185__C _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06347__S1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12523_ _01024_ net322 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12334__CLK net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12454_ _00955_ net252 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11548__A2 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11405_ u_cpu.rf_ram.memory\[26\]\[0\] _05683_ _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__A1 u_cpu.rf_ram.memory\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12385_ _00886_ net471 u_cpu.rf_ram.memory\[122\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11336_ u_cpu.rf_ram.memory\[88\]\[6\] _05626_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12484__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06975__A2 _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11267_ u_cpu.rf_ram.memory\[86\]\[5\] _05587_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13006_ _00066_ net528 u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _04717_ _04879_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11198_ _02976_ _05539_ _05546_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__A2 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10149_ _04690_ _04821_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09677__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout274_I net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09531__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07152__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout441_I net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09429__A1 _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__A1 u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07360_ _02900_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08101__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06311_ _01498_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07291_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _02757_ _02844_ _02846_ _02766_ _02847_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09030_ u_cpu.rf_ram.memory\[133\]\[2\] _04019_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06242_ _01513_ _01888_ _01521_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11701__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ _01499_ _01781_ _01794_ _01820_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08404__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__I1 u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06510__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09932_ _04622_ _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11851__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12977__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08168__A1 u_cpu.rf_ram.memory\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09863_ _04570_ _04571_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08610__I _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06718__A2 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10361__B _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07915__A1 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03853_ _03876_ _03882_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ u_arbiter.i_wb_cpu_rdt\[4\] _04512_ _04521_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08745_ u_cpu.rf_ram.memory\[72\]\[3\] _03836_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05957_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__C1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06026__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11475__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10278__A2 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08676_ _03794_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05888_ _01466_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06577__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07627_ _03103_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07558_ _02908_ _03056_ _03058_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06509_ _01941_ _02153_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08643__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07489_ u_cpu.rf_ram.memory\[18\]\[6\] _03003_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09228_ _04090_ _04140_ _04145_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ _03067_ _04013_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11211__I _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12170_ _00684_ net85 u_cpu.rf_ram.memory\[130\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11121_ u_cpu.rf_ram.memory\[108\]\[7\] _05488_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11052_ u_cpu.rf_ram.memory\[106\]\[7\] _05443_ _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07906__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10003_ _04655_ _04690_ _04692_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06040__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__A1 u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06590__B1 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11466__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10269__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11954_ _00476_ net37 u_cpu.rf_ram.memory\[55\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__S _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08331__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06568__S1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ _03453_ _05158_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06193__I0 u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11885_ _00407_ net87 u_cpu.rf_ram.memory\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06196__B _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10836_ _05320_ _05312_ _05321_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11724__CLK net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10767_ u_cpu.rf_ram.memory\[94\]\[4\] _05275_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12506_ _01007_ net172 u_cpu.rf_ram.memory\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10698_ _02467_ _05224_ _05225_ _04942_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06740__S1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12437_ _00938_ net246 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11874__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08398__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06215__I _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12368_ _00869_ net422 u_cpu.rf_ram.memory\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06799__I2 u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ _02913_ _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12299_ _00800_ net316 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08430__I _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout391_I net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout489_I net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06860_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07046__I _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ u_cpu.cpu.decode.op21 _01442_ _01460_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06791_ _01672_ _02432_ _01676_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06581__B1 _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__S0 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ _03673_ _03694_ _03701_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11457__A1 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06885__I _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08322__A1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__S1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ u_cpu.rf_ram.memory\[58\]\[4\] _03654_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08873__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07412_ _02909_ _02952_ _02953_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03537_ _03480_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _02878_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08625__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09822__A1 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07274_ _02832_ _02827_ _02783_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08605__I _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10356__B _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06731__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09013_ u_cpu.rf_ram.memory\[134\]\[5\] _04001_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06225_ _01692_ _01859_ _01872_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__13005__CLK net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08389__A1 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06156_ _01599_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10196__A1 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__A2 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10196__B2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06495__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06087_ _01637_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05964__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09915_ _04602_ _02646_ _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_113_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06247__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ _04518_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__A1 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _04486_ _04506_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06989_ _02495_ _02611_ _02464_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _03638_ _03820_ _03827_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11448__A1 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11747__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A1 u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06728__C _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ u_cpu.rf_ram.memory\[142\]\[1\] _03784_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10120__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11670_ _00192_ net464 u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10621_ _05171_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08616__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11897__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10552_ _05106_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06722__S1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _05084_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12222_ _00736_ net344 u_cpu.rf_ram.memory\[124\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06035__I _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09041__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10187__B2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06486__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12153_ _00667_ net77 u_cpu.rf_ram.memory\[132\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05874__I _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11104_ _05488_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07067__S _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12084_ _00598_ net63 u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11035_ _05443_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12522__CLK net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07355__A2 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__A1 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11439__A1 _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12986_ _00044_ net516 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07107__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12672__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__A1 _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11937_ _00459_ net38 u_cpu.rf_ram.memory\[57\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08855__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11868_ _00390_ net183 u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10819_ _03272_ _05308_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13028__CLK net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__A1 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout237_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08607__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11799_ _00321_ net18 u_cpu.rf_ram.memory\[74\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08425__I _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09280__A2 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06713__S1 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout404_I net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ _01510_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12052__CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09032__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10717__A3 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06477__S0 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09256__I _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _03181_ _03328_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09700_ u_cpu.rf_ram.memory\[115\]\[3\] _04451_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06912_ _02533_ _02550_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ _02524_ _02491_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08543__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ u_cpu.rf_ram.memory\[11\]\[3\] _04406_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06843_ _02462_ _02465_ _02483_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10350__A1 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06829__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09562_ _04364_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06774_ _01735_ _02415_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout52_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09099__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ u_cpu.rf_ram.memory\[56\]\[6\] _03686_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _04320_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10102__A1 _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10102__B2 _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08444_ _03644_ _03625_ _03645_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10653__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ u_cpu.rf_ram.memory\[60\]\[0\] _03598_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05959__I _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06609__A1 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10405__A2 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ _02484_ _02875_ _02869_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06704__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06208_ u_cpu.rf_ram.memory\[84\]\[1\] u_cpu.rf_ram.memory\[85\]\[1\] u_cpu.rf_ram.memory\[86\]\[1\]
+ u_cpu.rf_ram.memory\[87\]\[1\] _01855_ _01713_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05832__A2 _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07188_ _02701_ u_scanchain_local.module_data_in\[49\] _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10169__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06139_ u_cpu.rf_ram.memory\[0\]\[1\] u_cpu.rf_ram.memory\[1\]\[1\] u_cpu.rf_ram.memory\[2\]\[1\]
+ u_cpu.rf_ram.memory\[3\]\[1\] _01786_ _01553_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06468__S0 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12545__CLK net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05908__B _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07585__A2 _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout420 net421 net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout431 net434 net431 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout442 net443 net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout453 net460 net453 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout464 net468 net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout475 net476 net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08534__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout486 net489 net486 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout497 net498 net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09829_ u_arbiter.i_wb_cpu_rdt\[13\] _04546_ _04547_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10341__A1 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12840_ _01337_ net113 u_cpu.rf_ram.memory\[87\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12771_ _01268_ net129 u_cpu.rf_ram.memory\[108\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06848__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11722_ _00244_ net295 u_cpu.rf_ram.memory\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10644__A2 _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11653_ _00175_ net389 u_cpu.rf_ram.memory\[42\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net66 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05869__I _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A4 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout71 net74 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ u_cpu.rf_ram.memory\[109\]\[1\] _05161_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09798__B1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_11584_ _00106_ net410 u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _05120_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _05075_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09014__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10724__B _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12205_ _00719_ net298 u_cpu.rf_ram.memory\[126\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _04800_ _05035_ _05037_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07576__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08773__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12136_ _00650_ net62 u_cpu.rf_ram.memory\[134\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12067_ _00581_ net58 u_cpu.rf_ram.memory\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07328__A2 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _05399_ _05432_ _05434_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout187_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07324__I _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout354_I net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12969_ _00095_ net520 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10635__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06490_ u_cpu.rf_ram.memory\[44\]\[4\] u_cpu.rf_ram.memory\[45\]\[4\] u_cpu.rf_ram.memory\[46\]\[4\]
+ u_cpu.rf_ram.memory\[47\]\[4\] _01805_ _02030_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07500__A2 _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout521_I net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08160_ u_cpu.rf_ram.memory\[6\]\[2\] _03461_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10399__A1 _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02513_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06067__A2 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__A2 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ u_cpu.rf_ram.memory\[74\]\[2\] _03416_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ u_arbiter.i_wb_cpu_rdt\[7\] u_arbiter.i_wb_cpu_dbus_dat\[4\] _02652_ _02656_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05814__A2 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09005__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07567__A2 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06614__I1 u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08993_ _03729_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _03313_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07875_ u_cpu.rf_ram.memory\[4\]\[5\] _03263_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10323__A1 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09614_ u_cpu.rf_ram.memory\[8\]\[5\] _04393_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06826_ u_cpu.cpu.immdec.imm11_7\[0\] _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ u_cpu.rf_ram.memory\[120\]\[1\] _04354_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06757_ _02392_ _02394_ _02396_ _02398_ _01665_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08819__A2 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12098__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09476_ _04246_ _04309_ _04311_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06688_ _02055_ _02330_ _02058_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__A2 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08427_ u_cpu.rf_ram.memory\[5\]\[2\] _03632_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08358_ _03583_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07309_ _02852_ _02859_ _02862_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07255__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11051__A2 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ _03538_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10320_ _04721_ _04641_ _04709_ _04733_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05805__A2 _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11935__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _04714_ _04913_ _04854_ _04902_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07558__A2 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07409__I _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10182_ _04702_ _04704_ _04779_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06766__B1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10562__B2 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout250 net251 net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout261 net262 net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout272 net277 net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout283 net284 net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10314__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout294 net297 net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06469__B _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12823_ _01320_ net118 u_cpu.rf_ram.memory\[86\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12754_ _01251_ net116 u_cpu.rf_ram.memory\[107\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07494__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11705_ _00227_ net393 u_cpu.rf_ram.memory\[48\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12685_ _01182_ net170 u_cpu.rf_ram.memory\[101\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12710__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11636_ _00158_ net212 u_cpu.rf_ram.memory\[80\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09235__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07246__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11567_ _02585_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram_if.rtrig0 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07797__A2 _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08994__A1 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10518_ _05109_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11498_ u_cpu.rf_ram.memory\[98\]\[6\] _05734_ _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06651__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout102_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10449_ _05047_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08746__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10553__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12119_ _00633_ net283 u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06221__A2 _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ u_cpu.rf_ram.memory\[48\]\[0\] u_cpu.rf_ram.memory\[49\]\[0\] u_cpu.rf_ram.memory\[50\]\[0\]
+ u_cpu.rf_ram.memory\[51\]\[0\] _01636_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09534__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10305__A1 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__A1 u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07660_ u_cpu.rf_ram.memory\[46\]\[4\] _03122_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06604__S0 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06611_ _01580_ _02245_ _02254_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07591_ _03027_ _03071_ _03078_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__I0 u_cpu.rf_ram.memory\[120\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11808__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09330_ u_cpu.rf_ram.memory\[37\]\[5\] _04209_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10608__A2 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06542_ _02167_ _02186_ _01743_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ u_cpu.rf_ram.memory\[124\]\[4\] _04162_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06473_ _02006_ _02117_ _01728_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12390__CLK net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08212_ _03426_ _03483_ _03492_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout15_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09192_ _04095_ _04116_ _04123_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ u_cpu.rf_ram.memory\[75\]\[5\] _03446_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11033__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10092__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07788__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08985__A1 u_cpu.rf_ram.memory\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ u_cpu.rf_ram.memory\[77\]\[5\] _03401_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05799__A1 _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10792__A1 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ _02644_ _02635_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08976_ u_cpu.rf_ram.memory\[135\]\[0\] _03983_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ u_cpu.rf_ram.memory\[16\]\[3\] _03306_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10147__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__A1 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ _03228_ _03246_ _03255_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07712__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06809_ _02188_ _02450_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07789_ _02907_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12733__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09528_ _04167_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09459_ _04296_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12457__D _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__I0 u_cpu.rf_ram.memory\[92\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11272__A2 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11214__I _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10258__C _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12470_ _00971_ net490 u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05877__I2 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11421_ _05636_ _05683_ _05692_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07228__A1 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11024__A2 _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06752__B _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__A2 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08976__A1 u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11352_ _02616_ _02627_ _05647_ _03273_ _05644_ _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10783__A1 u_cpu.rf_ram.memory\[95\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10303_ _04716_ _04710_ _04958_ _04823_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11283_ u_cpu.rf_ram.memory\[111\]\[3\] _05599_ _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06451__A2 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08728__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13022_ _00084_ net534 u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06043__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ _04897_ _04673_ _04777_ _04748_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06203__A2 _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10165_ _04753_ _04729_ _04744_ _04820_ _04727_ _04835_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_117_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12263__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07951__A2 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10096_ _04764_ _04642_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10838__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08900__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12806_ _01303_ net111 u_cpu.rf_ram.memory\[85\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10998_ _05399_ _05420_ _05422_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07602__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07467__A1 u_cpu.rf_ram.memory\[81\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12737_ _01234_ net120 u_cpu.rf_ram.memory\[105\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11263__A2 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11124__I _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12668_ _01165_ net47 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09208__A2 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11619_ _00141_ net445 u_cpu.rf_ram.memory\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout317_I net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12599_ _01096_ net445 u_cpu.rf_ram.memory\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08433__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12606__CLK net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10526__B2 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _03848_ _03889_ _03892_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06888__I _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09264__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07942__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08761_ _03735_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05973_ _01511_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07712_ _03142_ _03155_ _03161_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08692_ u_cpu.rf_ram.memory\[141\]\[7\] _03794_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09695__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07643_ _03027_ _03107_ _03114_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07574_ _02884_ _03011_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07512__I _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09447__A2 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11780__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _04174_ _04194_ _04202_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07458__A1 u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06525_ u_cpu.rf_ram.memory\[88\]\[4\] u_cpu.rf_ram.memory\[89\]\[4\] u_cpu.rf_ram.memory\[90\]\[4\]
+ u_cpu.rf_ram.memory\[91\]\[4\] _01961_ _01674_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09244_ u_cpu.rf_ram.memory\[124\]\[0\] _04155_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06456_ u_cpu.rf_ram.memory\[132\]\[3\] u_cpu.rf_ram.memory\[133\]\[3\] u_cpu.rf_ram.memory\[134\]\[3\]
+ u_cpu.rf_ram.memory\[135\]\[3\] _02101_ _01754_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09175_ u_cpu.rf_ram.memory\[128\]\[6\] _04108_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06387_ _02023_ _02026_ _02029_ _02032_ _01613_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05967__I _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__A1 u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ u_cpu.rf_ram.memory\[76\]\[7\] _03428_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08057_ u_cpu.rf_ram.memory\[139\]\[7\] _03383_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07008_ _02630_ u_cpu.cpu.genblk3.csr.i_mtip _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10517__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09383__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08186__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06197__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06292__S1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08959_ _03930_ _03970_ _03973_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09135__A1 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11970_ _00492_ net38 u_cpu.rf_ram.memory\[53\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06339__I3 u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10921_ u_cpu.rf_ram.memory\[102\]\[6\] _05367_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06744__I0 u_cpu.rf_ram.memory\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06747__B _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10852_ _05332_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__I _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ u_cpu.rf_ram.memory\[95\]\[2\] _05287_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12522_ _01023_ net311 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06038__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12453_ _00954_ net252 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08949__A1 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _05681_ _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12629__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12384_ _00885_ net471 u_cpu.rf_ram.memory\[122\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _02944_ _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07621__A1 u_cpu.rf_ram.memory\[78\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06275__I2 u_cpu.rf_ram.memory\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11266_ _05562_ _05583_ _05590_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08177__A2 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13005_ _00065_ net527 u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10217_ _04876_ _04881_ _04883_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12779__CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ u_cpu.rf_ram.memory\[10\]\[4\] _05543_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11181__A1 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _04613_ _04691_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09126__A1 u_cpu.rf_ram.memory\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10079_ _04607_ _04690_ _04762_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12009__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09921__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout267_I net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09429__A2 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout434_I net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06310_ _01494_ _01946_ _01956_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07290_ _02757_ _02845_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06241_ u_cpu.rf_ram.memory\[24\]\[2\] u_cpu.rf_ram.memory\[25\]\[2\] u_cpu.rf_ram.memory\[26\]\[2\]
+ u_cpu.rf_ram.memory\[27\]\[2\] _01516_ _01774_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07860__A1 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09259__I _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06172_ _01795_ _01809_ _01819_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_8_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07612__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09931_ _04611_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09862_ u_arbiter.i_wb_cpu_rdt\[23\] _04495_ _04519_ u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout82_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__A3 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08813_ u_cpu.rf_ram.memory\[70\]\[3\] _03880_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _04496_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05956_ _01501_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_73_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08744_ _03739_ _03832_ _03837_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07128__B1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07128__C2 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07679__A1 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10868__I _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ _03794_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06026__S1 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11475__A2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05887_ _01509_ _01522_ _01527_ _01535_ _01490_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_96_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A2 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07626_ u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[4\] _02962_ _03085_
+ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ u_cpu.rf_ram.memory\[7\]\[0\] _03057_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06508_ u_cpu.rf_ram.memory\[108\]\[4\] u_cpu.rf_ram.memory\[109\]\[4\] u_cpu.rf_ram.memory\[110\]\[4\]
+ u_cpu.rf_ram.memory\[111\]\[4\] _02052_ _01827_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07488_ _02978_ _03000_ _03007_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09840__A2 _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06439_ _01555_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09227_ u_cpu.rf_ram.memory\[125\]\[2\] _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _04101_ _04086_ _04102_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ _03428_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07603__A1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ _04050_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _05484_ _05490_ _05498_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _05415_ _05445_ _05453_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11163__A1 _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10002_ _04655_ _04691_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05917__A1 _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10910__A1 u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__A1 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__A2 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06590__B2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11466__A2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11953_ _00475_ net25 u_cpu.rf_ram.memory\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08331__A2 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ _05328_ _05352_ _05361_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08248__I _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11884_ _00406_ net86 u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10835_ u_cpu.rf_ram.memory\[28\]\[3\] _05318_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06893__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06991__I _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08095__A1 _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10766_ _05209_ _05271_ _05277_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12451__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09831__A2 _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12505_ _01006_ net186 u_cpu.rf_ram.memory\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10697_ u_cpu.cpu.immdec.imm11_7\[1\] _04674_ _05224_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12436_ _00937_ net246 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10729__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09595__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08398__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12367_ _00868_ net422 u_cpu.rf_ram.memory\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09807__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11318_ _05618_ _05620_ _05622_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06799__I3 u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12298_ _00799_ net315 u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09347__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11249_ u_cpu.rf_ram.memory\[110\]\[6\] _05575_ _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11154__A1 u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09898__A2 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout384_I net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10901__A1 u_cpu.rf_ram.memory\[101\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ u_cpu.cpu.genblk3.csr.o_new_irq _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06790_ u_cpu.rf_ram.memory\[88\]\[7\] u_cpu.rf_ram.memory\[89\]\[7\] u_cpu.rf_ram.memory\[90\]\[7\]
+ u_cpu.rf_ram.memory\[91\]\[7\] _01673_ _01674_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09542__I _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10688__I _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11457__A2 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08322__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08460_ _03573_ _03650_ _03656_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07411_ u_cpu.rf_ram.memory\[82\]\[7\] _02900_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11209__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08391_ _03581_ _03598_ _03607_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06884__A2 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07342_ _02890_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09822__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07273_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12944__CLK net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09012_ _03748_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _01861_ _01866_ _01869_ _01871_ _01740_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06406__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08389__A2 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09586__A1 _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06155_ u_cpu.rf_ram.memory\[40\]\[1\] u_cpu.rf_ram.memory\[41\]\[1\] u_cpu.rf_ram.memory\[42\]\[1\]
+ u_cpu.rf_ram.memory\[43\]\[1\] _01569_ _01601_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11393__A1 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10196__A2 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06086_ _01710_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06495__S1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09914_ _04605_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09889__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08010__A1 _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06247__S1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09845_ _04494_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12324__CLK net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__I2 u_cpu.rf_ram.memory\[106\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09776_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _02649_ _02651_ _04487_ _04506_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06572__A1 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06988_ u_cpu.cpu.bufreg.lsb\[0\] _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05980__I _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08727_ u_cpu.rf_ram.memory\[13\]\[4\] _03824_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10598__I _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11448__A2 _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05939_ _01582_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08313__A2 _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _03730_ _03783_ _03785_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A2 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ _03018_ _03089_ _03092_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08589_ _03738_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10620_ _05171_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08077__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10959__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07700__I _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09813__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _05129_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10266__C _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06316__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10482_ u_cpu.cpu.bufreg.i_sh_signed u_arbiter.i_wb_cpu_dbus_adr\[31\] _02874_ _05085_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09577__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12221_ _00735_ net348 u_cpu.rf_ram.memory\[124\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__A2 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12152_ _00666_ net77 u_cpu.rf_ram.memory\[132\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06486__S1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10282__B _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11103_ _03152_ _05455_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09329__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12083_ _00597_ net63 u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11136__A1 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11034_ _03101_ _05374_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06051__I _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08001__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08552__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06402__I2 u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__A1 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05890__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07083__S _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11439__A2 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12985_ _00043_ net516 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09501__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11936_ _00458_ net67 u_cpu.rf_ram.memory\[57\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10111__A2 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _00389_ net183 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11841__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12967__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08068__A1 u_cpu.rf_ram.memory\[77\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10818_ _02715_ _05307_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11798_ _00320_ net15 u_cpu.rf_ram.memory\[74\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout132_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10749_ u_cpu.rf_ram.memory\[97\]\[5\] _05263_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06174__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__A2 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09568__A1 u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12419_ _00920_ net248 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__A2 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11375__A1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08441__I _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08240__A1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06477__S1 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12347__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08791__A2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07960_ _03327_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11127__A1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ _02536_ _02537_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07891_ _03272_ _03279_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09630_ _04070_ _04402_ _04407_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06842_ _02462_ _02482_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12497__CLK net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10350__A2 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09272__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06773_ u_cpu.rf_ram.memory\[108\]\[7\] u_cpu.rf_ram.memory\[109\]\[7\] u_cpu.rf_ram.memory\[110\]\[7\]
+ u_cpu.rf_ram.memory\[111\]\[7\] _02052_ _01506_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09561_ _04364_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08512_ _03675_ _03683_ _03690_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09492_ _02890_ _03130_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06306__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout45_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10102__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08443_ u_cpu.rf_ram.memory\[5\]\[6\] _03632_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _03596_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ _02870_ _02872_ _02873_ _02874_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06165__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07256_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] u_cpu.cpu.ctrl.o_ibus_adr\[23\] _02810_ _02818_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_30_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06207_ _01502_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09559__A1 _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07187_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _02757_ _02760_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10169__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11366__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05975__I _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ _01549_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08231__A1 _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06468__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A2 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ _01697_ _01703_ _01709_ _01716_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11118__A1 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__I2 u_cpu.rf_ram.memory\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout410 net412 net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06793__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout421 net427 net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout432 net434 net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11714__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout443 net448 net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout454 net455 net454 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout465 net468 net465 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__A2 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout476 net484 net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout487 net489 net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09828_ _04518_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout498 net503 net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10341__A2 _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09759_ _03291_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11864__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10121__I _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12770_ _01267_ net138 u_cpu.rf_ram.memory\[108\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09910__I _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _00243_ net387 u_cpu.rf_ram.memory\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06848__A2 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11652_ _00174_ net389 u_cpu.rf_ram.memory\[42\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06474__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout61 net65 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_10603_ _04800_ _05160_ _05162_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09798__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout72 net74 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09798__B2 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout83 net93 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11583_ _00105_ net410 u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_31_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06046__I _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _05116_ _05118_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08470__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10465_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _05072_
+ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05885__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07078__S _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12204_ _00718_ net296 u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10396_ u_cpu.rf_ram.memory\[31\]\[0\] _05036_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06084__I0 u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09970__A1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12135_ _00649_ net43 u_cpu.rf_ram.memory\[134\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08773__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11109__A1 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10580__A2 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12066_ _00580_ net15 u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ u_cpu.rf_ram.memory\[105\]\[0\] _05433_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12968_ _00094_ net520 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10096__A1 _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11919_ _00441_ net221 u_cpu.rf_ram.memory\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10966__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout347_I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12899_ _01396_ net437 u_cpu.rf_ram.memory\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06395__S0 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__A1 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10399__A2 _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07110_ _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _03409_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A1 u_cpu.rf_ram.memory\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07041_ _02655_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09267__I _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06224__B1 _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ _03943_ _03983_ _03992_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07943_ _03215_ _03314_ _03317_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11887__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__A1 u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08516__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07874_ _02934_ _03259_ _03266_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10323__A2 _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07515__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04075_ _04389_ _04396_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06825_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ _04332_ _04353_ _04355_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06756_ _01538_ _02397_ _01663_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10087__A1 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09475_ u_cpu.rf_ram.memory\[35\]\[0\] _04310_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06687_ u_cpu.rf_ram.memory\[104\]\[6\] u_cpu.rf_ram.memory\[105\]\[6\] u_cpu.rf_ram.memory\[106\]\[6\]
+ u_cpu.rf_ram.memory\[107\]\[6\] _02056_ _01624_ _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_19_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08426_ _03623_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _03568_ _03584_ _03587_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12512__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ _02860_ _02861_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__A1 u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08288_ _03498_ _03539_ _03542_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ _02800_ _02802_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11339__A1 u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10250_ u_arbiter.i_wb_cpu_rdt\[29\] u_arbiter.i_wb_cpu_rdt\[13\] _04773_ _04913_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08204__A1 _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _04790_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06766__B2 _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout240 net243 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout251 net256 net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout262 net267 net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08507__A2 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout273 net275 net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11511__A1 _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout284 net290 net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout295 net297 net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07191__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12822_ _01319_ net111 u_cpu.rf_ram.memory\[86\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12753_ _01250_ net116 u_cpu.rf_ram.memory\[107\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10873__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11704_ _00226_ net296 u_cpu.rf_ram.memory\[48\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12684_ _01181_ net170 u_cpu.rf_ram.memory\[101\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08691__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11635_ _00157_ net208 u_cpu.rf_ram.memory\[80\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12192__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06129__S0 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11566_ _05779_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _03270_ _02865_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08994__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11497_ _03640_ _05731_ _05738_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10448_ _05065_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10379_ _04805_ _05023_ _05026_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06757__A1 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06301__S0 _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12118_ _00632_ net265 u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout297_I net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12049_ _00563_ net33 u_cpu.rf_ram.memory\[73\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06509__A1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11502__A1 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10305__A2 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09171__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout464_I net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06604__S1 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06610_ _02247_ _02249_ _02251_ _02253_ _02072_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07590_ u_cpu.rf_ram.memory\[80\]\[5\] _03074_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10069__A1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06541_ _01958_ _02176_ _02185_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06368__S0 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12535__CLK net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06472_ u_cpu.rf_ram.memory\[16\]\[4\] u_cpu.rf_ram.memory\[17\]\[4\] u_cpu.rf_ram.memory\[18\]\[4\]
+ u_cpu.rf_ram.memory\[19\]\[4\] _02007_ _01518_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10864__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ _04167_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07485__A2 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ u_cpu.rf_ram.memory\[67\]\[7\] _03481_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09191_ u_cpu.rf_ram.memory\[127\]\[4\] _04120_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11569__A1 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _03420_ _03442_ _03449_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10241__A1 _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ _03344_ _03397_ _03404_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10092__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08985__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06996__A1 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__A2 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10792__A2 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07024_ _02612_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09934__A1 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10544__A2 _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ _03981_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ _03217_ _03302_ _03307_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07857_ u_cpu.rf_ram.memory\[50\]\[7\] _03244_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06808_ u_cpu.rf_ram.memory\[128\]\[7\] u_cpu.rf_ram.memory\[129\]\[7\] u_cpu.rf_ram.memory\[130\]\[7\]
+ u_cpu.rf_ram.memory\[131\]\[7\] _01764_ _01765_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07788_ _03150_ _03200_ _03209_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06920__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ _04342_ _04334_ _04343_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06739_ _02374_ _02376_ _02378_ _02380_ _01717_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10855__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07476__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09458_ _04251_ _04297_ _04300_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08673__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09870__B1 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08409_ _03579_ _03610_ _03618_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09389_ u_cpu.rf_ram.memory\[91\]\[1\] _04249_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11420_ u_cpu.rf_ram.memory\[26\]\[7\] _05681_ _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07228__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08804__I _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10232__A1 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11351_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11230__I _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10783__A2 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10302_ _04747_ _04628_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06324__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _05557_ _05595_ _05600_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06451__A3 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08728__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13021_ _00083_ net534 u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10233_ _04636_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06739__A1 _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10164_ _04824_ _04834_ _04836_ _04689_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_121_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10290__B _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10095_ _04672_ _04777_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07164__A1 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06911__A1 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12805_ _01302_ net103 u_cpu.rf_ram.memory\[85\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10997_ u_cpu.rf_ram.memory\[79\]\[0\] _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12736_ _01233_ net148 u_cpu.rf_ram.memory\[105\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07467__A2 _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08664__A1 u_cpu.rf_ram.memory\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12667_ _01164_ net175 u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11618_ _00140_ net498 u_cpu.rf_ram.memory\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07219__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12598_ _01095_ net441 u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06427__B1 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10223__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout212_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11549_ _05765_ _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10774__A2 _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08719__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10526__A2 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ _03843_ _03845_ _03847_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05972_ _01615_ _01620_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07711_ u_cpu.rf_ram.memory\[44\]\[3\] _03159_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08691_ _03752_ _03796_ _03804_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07155__A1 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06202__I0 u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07642_ u_cpu.rf_ram.memory\[42\]\[5\] _03110_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06753__I1 u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ _02952_ _03057_ _03066_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11315__I _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09312_ u_cpu.rf_ram.memory\[38\]\[6\] _04197_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06524_ _01693_ _02168_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07014__B _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06409__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ _04153_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06455_ _01746_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08407__A1 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06386_ _01915_ _02031_ _01807_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09174_ _04097_ _04105_ _04112_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06572__C _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06269__I0 u_cpu.rf_ram.memory\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ _03424_ _03430_ _03438_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06513__S0 _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10765__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06144__I _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ _03350_ _03385_ _03393_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07007_ _02629_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10517__A2 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09383__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11190__A2 _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08958_ u_cpu.rf_ram.memory\[136\]\[1\] _03971_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09135__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _02885_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _03296_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07146__A1 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08889_ u_cpu.rf_ram.memory\[39\]\[0\] _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10920_ _05324_ _05364_ _05371_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06744__I1 u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10851_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _05331_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07161__A4 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10782_ _05282_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12521_ _01022_ net322 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06121__A2 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12452_ _00953_ net474 u_cpu.rf_ram.memory\[113\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10205__A1 _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11403_ _05681_ _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08949__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12383_ _00884_ net471 u_cpu.rf_ram.memory\[122\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09071__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06504__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11334_ _05632_ _05621_ _05633_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ u_cpu.rf_ram.memory\[86\]\[4\] _05587_ _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10508__A2 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05893__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13004_ _00064_ net527 u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10216_ u_cpu.cpu.immdec.imm30_25\[0\] _04882_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11196_ _02974_ _05539_ _05545_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06432__I0 u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11181__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _02708_ _04820_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11948__CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A2 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07137__A1 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10078_ _04692_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07688__A2 _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout162_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12719_ _01216_ net155 u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout427_I net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06673__B _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ _01500_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07860__A2 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06171_ _01811_ _01814_ _01816_ _01818_ _01642_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09062__A1 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10747__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _03275_ u_arbiter.i_wb_cpu_rdt\[0\] _04621_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09275__I _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _04521_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11172__A2 _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _03850_ _03876_ _03881_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07009__B _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _04490_ _04517_ _04519_ _04520_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout75_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05926__A2 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09117__A2 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12873__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08743_ u_cpu.rf_ram.memory\[72\]\[2\] _03836_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05955_ _01537_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07679__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08876__A1 _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _03131_ _03370_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05886_ _01528_ _01531_ _01534_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07625_ _03101_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12103__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08628__A1 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07556_ _03055_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06507_ _01937_ _02151_ _01596_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ u_cpu.rf_ram.memory\[18\]\[5\] _03003_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10986__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _04139_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06438_ u_cpu.rf_ram.memory\[84\]\[3\] u_cpu.rf_ram.memory\[85\]\[3\] u_cpu.rf_ram.memory\[86\]\[3\]
+ u_cpu.rf_ram.memory\[87\]\[3\] _01855_ _02083_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12253__CLK net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09157_ u_cpu.rf_ram.memory\[22\]\[7\] _04084_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09053__A1 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06369_ _01785_ _02014_ _01902_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10199__B1 _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10738__A2 _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08108_ _03395_ _03153_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07603__A2 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _03998_ _04051_ _04054_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08800__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06257__I3 u_cpu.rf_ram.memory\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ _03196_ _03370_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11050_ u_cpu.rf_ram.memory\[106\]\[6\] _05448_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11163__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10001_ _04663_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__I1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09913__I _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06590__A2 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11952_ _00474_ net25 u_cpu.rf_ram.memory\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10674__A1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10903_ u_cpu.rf_ram.memory\[101\]\[7\] _05350_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11883_ _00405_ net86 u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06342__A2 _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08619__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10834_ _05208_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06049__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12926__D _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ u_cpu.rf_ram.memory\[94\]\[3\] _05275_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08095__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10977__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05888__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12504_ _01005_ net186 u_cpu.rf_ram.memory\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A2 _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10696_ _03278_ _05223_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12435_ _00936_ net236 u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11620__CLK net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10729__A2 _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12366_ _00867_ net422 u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11317_ u_cpu.rf_ram.memory\[88\]\[0\] _05621_ _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12297_ _00798_ net255 u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09347__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11770__CLK net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11248_ _05564_ _05572_ _05579_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__I _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11179_ _05482_ _05527_ _05534_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05908__A2 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__I _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout377_I net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06668__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08858__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07343__I _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__A1 _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__C _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ _02951_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12276__CLK net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ u_cpu.rf_ram.memory\[60\]\[7\] _03596_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07341_ _02884_ _02889_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11090__A1 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__B1 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08174__I _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ u_scanchain_local.module_data_in\[64\] _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07833__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05844__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _04005_ _03995_ _04006_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06223_ _01735_ _01870_ _01738_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09035__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06154_ _01589_ _01800_ _01801_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09586__A2 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07597__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11393__A2 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ _01730_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07518__I _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _04604_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__A1 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09844_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _04557_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08010__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _04487_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__I3 u_cpu.rf_ram.memory\[107\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06987_ u_cpu.cpu.bufreg.lsb\[1\] _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08726_ _03635_ _03820_ _03826_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10105__B1 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05938_ u_cpu.rf_ram.memory\[36\]\[0\] u_cpu.rf_ram.memory\[37\]\[0\] u_cpu.rf_ram.memory\[38\]\[0\]
+ u_cpu.rf_ram.memory\[39\]\[0\] _01584_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12619__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10656__A1 _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ u_cpu.rf_ram.memory\[142\]\[0\] _03784_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05869_ _01517_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07608_ u_cpu.rf_ram.memory\[78\]\[1\] _03090_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _02918_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10408__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ u_cpu.rf_ram.memory\[1\]\[3\] _03043_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08077__A2 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09274__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11503__I _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12769__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10550_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _05123_ _05125_ _02769_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07824__A2 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09209_ u_cpu.rf_ram.memory\[126\]\[3\] _04132_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__I _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09026__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10481_ _02856_ _02858_ _05083_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09908__I _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12220_ _00734_ net350 u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11793__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09577__A2 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12151_ _00665_ net52 u_cpu.rf_ram.memory\[132\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06260__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _05486_ _05471_ _05487_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06332__I _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12082_ _00596_ net222 u_cpu.rf_ram.memory\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12149__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11136__A2 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _05417_ _05433_ _05442_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08001__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__I _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07760__A1 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12984_ _00042_ net513 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12299__CLK net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09501__A2 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11935_ _00457_ net69 u_cpu.rf_ram.memory\[57\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11866_ _00388_ net106 u_cpu.rf_ram.memory\[64\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _02699_ _02632_ _02702_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08068__A2 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A1 u_cpu.rf_ram.memory\[124\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11797_ _00319_ net15 u_cpu.rf_ram.memory\[74\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11072__A1 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _05212_ _05259_ _05266_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07815__A2 _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06174__S1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05826__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout125_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09017__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10679_ _02931_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12418_ _00919_ net248 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11375__A2 _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12349_ _00850_ net472 u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08240__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout494_I net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11127__A2 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06910_ u_cpu.cpu.bufreg.lsb\[0\] _02530_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07890_ _03273_ u_cpu.cpu.state.stage_two_req _03278_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_25_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07051__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09740__A2 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ _02466_ _02479_ _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07751__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _03355_ _03453_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06772_ _01589_ _02413_ _01596_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10638__A1 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08511_ u_cpu.rf_ram.memory\[56\]\[5\] _03686_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09491_ _04264_ _04310_ _04319_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11666__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06306__A2 _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _03643_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12911__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout38_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03596_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11323__I _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10367__C _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07324_ _02864_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06165__S1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10810__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ _02701_ u_scanchain_local.module_data_in\[61\] _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09008__A1 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06206_ _01852_ _01853_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07186_ _02758_ _02753_ _02759_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10169__A3 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ _01512_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10574__B1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _01489_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout400 net407 net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout411 net412 net411 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11118__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout422 net426 net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07990__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout433 net434 net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout444 net448 net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05991__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout455 net459 net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout466 net467 net466 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12441__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07042__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09827_ _04494_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout477 net480 net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout488 net489 net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout499 net503 net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06545__A2 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _03282_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _03749_ _03808_ _03815_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04444_ _04429_ _04445_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12591__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11720_ _00242_ net295 u_cpu.rf_ram.memory\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11651_ _00173_ net389 u_cpu.rf_ram.memory\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout40 net41 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net54 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10602_ u_cpu.rf_ram.memory\[109\]\[0\] _05161_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout62 net65 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_54_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11582_ _00104_ net410 u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout73 net74 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_141_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout84 net88 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10801__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10533_ _05119_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__A2 _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10464_ _05074_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12203_ _00717_ net296 u_cpu.rf_ram.memory\[126\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10395_ _05034_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10565__B1 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06062__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12134_ _00648_ net52 u_cpu.rf_ram.memory\[134\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06084__I1 u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09970__A2 _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11109__A2 _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06997__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12065_ _00579_ net10 u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11016_ _05431_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09722__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11689__CLK net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07733__A1 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12934__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12967_ _00093_ net519 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11918_ _00440_ net220 u_cpu.rf_ram.memory\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11293__A1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10096__A2 _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12898_ _01395_ net438 u_cpu.rf_ram.memory\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11849_ _00371_ net98 u_cpu.rf_ram.memory\[66\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout242_I net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09238__A1 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11143__I _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10187__C _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A1 _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10982__I _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12314__CLK net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout507_I net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08461__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ u_arbiter.i_wb_cpu_rdt\[6\] u_arbiter.i_wb_cpu_dbus_dat\[3\] _02652_ _02655_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10556__B1 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ u_cpu.rf_ram.memory\[135\]\[7\] _03981_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06614__I3 u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ u_cpu.rf_ram.memory\[17\]\[1\] _03315_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10423__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09283__I _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__A2 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07873_ u_cpu.rf_ram.memory\[4\]\[4\] _03263_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07724__A1 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ u_cpu.rf_ram.memory\[8\]\[4\] _04393_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11520__A2 _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06824_ _02463_ u_cpu.cpu.bufreg.i_sh_signed _02464_ _01444_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09543_ u_cpu.rf_ram.memory\[120\]\[0\] _04354_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06755_ u_cpu.rf_ram.memory\[44\]\[7\] u_cpu.rf_ram.memory\[45\]\[7\] u_cpu.rf_ram.memory\[46\]\[7\]
+ u_cpu.rf_ram.memory\[47\]\[7\] _01661_ _02030_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06856__B _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11284__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ _04308_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06686_ _01941_ _02328_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07531__I _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08425_ _03630_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06147__I _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08356_ u_cpu.rf_ram.memory\[61\]\[1\] _03585_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ u_cpu.cpu.state.stage_two_req _02529_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10892__I _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08287_ u_cpu.rf_ram.memory\[29\]\[1\] _03540_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05986__I _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07238_ _02800_ _02802_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11339__A2 _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07169_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _02740_ _02713_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08204__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10011__A2 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _02708_ _04849_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06766__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12957__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout230 net231 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout241 net243 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__A2 _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout252 net254 net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout263 net266 net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout274 net275 net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07715__A1 u_cpu.rf_ram.memory\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06518__A2 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout285 net289 net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout296 net297 net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10132__I _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11981__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12821_ _01318_ net101 u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 u_cpu.rf_ram.memory\[92\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12752_ _01249_ net145 u_cpu.rf_ram.memory\[107\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08140__A1 _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11703_ _00225_ net387 u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12683_ _01180_ net46 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08691__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11027__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _00156_ net212 u_cpu.rf_ram.memory\[80\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06057__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06129__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11565_ _02585_ _02587_ u_cpu.rf_ram.rdata\[7\] _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08443__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__A1 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07089__S _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06454__A1 _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10516_ _05107_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12487__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11496_ u_cpu.rf_ram.memory\[98\]\[5\] _05734_ _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10447_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _05060_
+ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06006__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06206__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ u_cpu.rf_ram.memory\[32\]\[1\] _05024_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07954__A1 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06301__S1 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12117_ _00631_ net265 u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ _00562_ net33 u_cpu.rf_ram.memory\[73\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout192_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07706__A1 u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11502__A2 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06065__S0 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__A1 _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02178_ _02180_ _02182_ _02184_ _01982_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__S1 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _01890_ _02115_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08682__A2 _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08210_ _03424_ _03483_ _03491_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11018__A1 _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06693__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09190_ _04093_ _04116_ _04122_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11704__CLK net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ u_cpu.rf_ram.memory\[75\]\[4\] _03446_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__I _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08072_ u_cpu.rf_ram.memory\[77\]\[4\] _03401_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10241__A2 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06996__A2 _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07023_ _02629_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11854__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10529__B1 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08198__A1 u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08910__I _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06599__I2 u_cpu.rf_ram.memory\[106\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08974_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ u_cpu.rf_ram.memory\[16\]\[2\] _03306_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ _03226_ _03246_ _03254_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08370__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06807_ _02429_ _02448_ _01475_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10887__I _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ u_cpu.rf_ram.memory\[43\]\[7\] _03198_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06920__A2 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11257__A1 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ u_cpu.rf_ram.memory\[117\]\[3\] _04340_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06738_ _02006_ _02379_ _01728_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09457_ u_cpu.rf_ram.memory\[92\]\[1\] _04298_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06669_ _02305_ _02307_ _02309_ _02311_ _01665_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09870__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08673__A2 _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11009__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ u_cpu.rf_ram.memory\[19\]\[6\] _03613_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09388_ _04157_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08339_ _03343_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11350_ _02504_ _05641_ _05646_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10301_ _04956_ _04948_ _04957_ _04758_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11281_ u_cpu.rf_ram.memory\[111\]\[2\] _05599_ _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08189__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13020_ _00082_ net534 u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09916__I _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10232_ _04895_ _04896_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07936__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__S0 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _04608_ _04781_ _04777_ _04835_ _04653_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07436__I _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09689__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ _04732_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06047__S0 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11496__A1 u_cpu.rf_ram.memory\[98\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__I _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11248__A1 _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12804_ _01301_ net100 u_cpu.rf_ram.memory\[85\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10996_ _05419_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12735_ _01232_ net148 u_cpu.rf_ram.memory\[105\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09861__A1 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08664__A2 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12666_ _01163_ net177 u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11617_ _00139_ net504 u_cpu.rf_ram.memory\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__A1 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12597_ _01094_ net441 u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10223__A2 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11548_ _03627_ _05766_ _05769_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06978__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10037__I _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout205_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11479_ _02980_ _05719_ _05727_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07927__A1 u_cpu.rf_ram.memory\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06250__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05971_ u_cpu.rf_ram.memory\[60\]\[0\] u_cpu.rf_ram.memory\[61\]\[0\] u_cpu.rf_ram.memory\[62\]\[0\]
+ u_cpu.rf_ram.memory\[63\]\[0\] _01617_ _01619_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07710_ _03139_ _03155_ _03160_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11487__A1 u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ u_cpu.rf_ram.memory\[141\]\[6\] _03799_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06202__I1 u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07641_ _03025_ _03106_ _03113_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11239__A1 _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07572_ u_cpu.rf_ram.memory\[7\]\[7\] _03055_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08104__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12652__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09311_ _04171_ _04194_ _04201_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06523_ u_cpu.rf_ram.memory\[92\]\[4\] u_cpu.rf_ram.memory\[93\]\[4\] u_cpu.rf_ram.memory\[94\]\[4\]
+ u_cpu.rf_ram.memory\[95\]\[4\] _02075_ _01847_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06666__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ _04153_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06454_ _01469_ _02099_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout20_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13008__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09173_ u_cpu.rf_ram.memory\[128\]\[5\] _04108_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09604__A1 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06385_ u_cpu.rf_ram.memory\[44\]\[3\] u_cpu.rf_ram.memory\[45\]\[3\] u_cpu.rf_ram.memory\[46\]\[3\]
+ u_cpu.rf_ram.memory\[47\]\[3\] _01805_ _02030_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08407__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06418__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08124_ u_cpu.rf_ram.memory\[76\]\[6\] _03433_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11411__A1 _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10214__A2 _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09080__A2 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06969__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06513__S1 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08055_ u_cpu.rf_ram.memory\[139\]\[6\] _03388_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12032__CLK net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07006_ _02628_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06277__S0 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08591__A1 u_cpu.rf_ram.memory\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08957_ _03925_ _03970_ _03972_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12182__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07908_ _02885_ _03295_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08888_ _03926_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07146__A2 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ _02891_ _03168_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10850_ _05330_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09509_ _04262_ _04322_ _04330_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _05202_ _05283_ _05286_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12520_ _01021_ net311 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12451_ _00952_ net481 u_cpu.rf_ram.memory\[113\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11402_ _05310_ _03102_ _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10285__C _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__A1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10205__A2 _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12382_ _00883_ net472 u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06335__I _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A2 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06504__S1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ u_cpu.rf_ram.memory\[88\]\[5\] _05626_ _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11264_ _05560_ _05583_ _05589_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13003_ _00063_ net527 u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12525__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _03278_ _04879_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11195_ u_cpu.rf_ram.memory\[10\]\[3\] _05543_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06070__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__I1 u_cpu.rf_ram.memory\[89\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _04818_ _04803_ _04819_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10077_ _04649_ _04666_ _04631_ _04608_ _04684_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_47_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12659__D _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__I2 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06896__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10979_ _05208_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06648__A1 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12718_ _01215_ net155 u_cpu.rf_ram.memory\[99\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06499__I1 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout322_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12649_ _01146_ net144 u_cpu.rf_ram.memory\[95\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11151__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12055__CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _01634_ _01817_ _01640_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__C _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09062__A2 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06259__S0 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09860_ _04568_ _04569_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07376__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ u_cpu.rf_ram.memory\[70\]\[2\] _03880_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09791_ _04518_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _03831_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05954_ _01599_ _01602_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout68_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ _03755_ _03784_ _03793_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05885_ _01533_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11326__I _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06726__I2 u_cpu.rf_ram.memory\[142\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06887__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07624_ _02889_ _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_78_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07555_ _03055_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08628__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06506_ u_cpu.rf_ram.memory\[96\]\[4\] u_cpu.rf_ram.memory\[97\]\[4\] u_cpu.rf_ram.memory\[98\]\[4\]
+ u_cpu.rf_ram.memory\[99\]\[4\] _01938_ _01824_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07486_ _02976_ _02999_ _03006_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _04088_ _04140_ _04143_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06437_ _01562_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09156_ _03754_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06368_ u_cpu.rf_ram.memory\[0\]\[3\] u_cpu.rf_ram.memory\[1\]\[3\] u_cpu.rf_ram.memory\[2\]\[3\]
+ u_cpu.rf_ram.memory\[3\]\[3\] _01786_ _01900_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10199__A1 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09053__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10199__B2 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08107_ _03426_ _03411_ _03427_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09087_ u_cpu.rf_ram.memory\[130\]\[1\] _04052_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06299_ _01936_ _01940_ _01943_ _01945_ _01832_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08800__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06811__A1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ _03353_ _03373_ _03382_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10000_ _04627_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09989_ _04596_ u_arbiter.i_wb_cpu_rdt\[4\] _04678_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_40_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06670__S0 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__A1 _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11951_ _00473_ net25 u_cpu.rf_ram.memory\[55\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10902_ _05326_ _05352_ _05360_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10674__A2 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11882_ _00404_ net167 u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _05317_ _05312_ _05319_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12078__CLK net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10764_ _05205_ _05271_ _05276_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12503_ _01004_ net490 u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10695_ _02618_ _02873_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12434_ _00935_ net235 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12365_ _00866_ net422 u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11316_ _05619_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06802__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11915__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12296_ _00797_ net314 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ u_cpu.rf_ram.memory\[110\]\[5\] _05575_ _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10315__I _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11178_ u_cpu.rf_ram.memory\[59\]\[5\] _05530_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10362__A1 _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _04801_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06661__S0 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08307__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout272_I net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08858__A2 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11146__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__A2 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05916__I0 u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10985__I _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout537_I net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06684__B _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07340_ _01591_ _02888_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07271_ _02827_ _02829_ _02830_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07294__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11090__A2 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__B2 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09010_ u_cpu.rf_ram.memory\[134\]\[4\] _04001_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06222_ u_cpu.rf_ram.memory\[76\]\[1\] u_cpu.rf_ram.memory\[77\]\[1\] u_cpu.rf_ram.memory\[78\]\[1\]
+ u_cpu.rf_ram.memory\[79\]\[1\] _01515_ _01736_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05844__A2 _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A2 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06153_ _01532_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11595__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10050__B1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__A1 _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06084_ u_cpu.rf_ram.memory\[72\]\[0\] u_cpu.rf_ram.memory\[73\]\[0\] u_cpu.rf_ram.memory\[74\]\[0\]
+ u_cpu.rf_ram.memory\[75\]\[0\] _01731_ _01732_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09912_ _04603_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_63_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08546__A1 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09843_ _04496_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10353__A1 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06652__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12990__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09774_ _04504_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06986_ net3 _02609_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08725_ u_cpu.rf_ram.memory\[13\]\[3\] _03824_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05937_ _01585_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10105__A1 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A2 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11056__I _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10105__B2 _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10656__A2 _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06404__S0 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _03782_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05868_ _01505_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12220__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07607_ _03010_ _03089_ _03091_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08587_ _03736_ _03732_ _03737_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05799_ _01448_ u_cpu.cpu.decode.op26 _01449_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05989__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07538_ _02921_ _03039_ _03044_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ u_cpu.rf_ram.memory\[81\]\[6\] _02991_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05835__A2 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09208_ _04090_ _04128_ _04133_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10480_ _02856_ _02858_ _02874_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11938__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09026__A2 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09139_ _04088_ _04085_ _04089_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07588__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12150_ _00664_ net53 u_cpu.rf_ram.memory\[132\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11101_ u_cpu.rf_ram.memory\[83\]\[7\] _05469_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12081_ _00595_ net222 u_cpu.rf_ram.memory\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06260__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10135__I _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08537__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11032_ u_cpu.rf_ram.memory\[105\]\[7\] _05431_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06643__S0 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12983_ _00041_ net513 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12002__D _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10647__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11934_ _00456_ net71 u_cpu.rf_ram.memory\[57\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _00387_ net105 u_cpu.rf_ram.memory\[64\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12713__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05899__I _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10816_ _04923_ _05306_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11796_ _00318_ net34 u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11072__A2 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10747_ u_cpu.rf_ram.memory\[97\]\[4\] _05263_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05826__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10678_ _05209_ _05198_ _05210_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09017__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12863__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07028__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12417_ _00918_ net247 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout118_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07579__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12348_ _00849_ net452 u_cpu.rf_ram.memory\[118\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12279_ _00780_ net313 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08528__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout487_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10335__A1 _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _02480_ u_cpu.cpu.alu.add_cy_r _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07051__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06634__S0 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__I _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12243__CLK net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ u_cpu.rf_ram.memory\[96\]\[7\] u_cpu.rf_ram.memory\[97\]\[7\] u_cpu.rf_ram.memory\[98\]\[7\]
+ u_cpu.rf_ram.memory\[99\]\[7\] _01590_ _01593_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08510_ _03673_ _03682_ _03689_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10638__A2 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09490_ u_cpu.rf_ram.memory\[35\]\[7\] _04308_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07503__A2 _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08700__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08441_ _02944_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08372_ _03152_ _03595_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07323_ _02558_ _02463_ _02578_ _02557_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_108_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ _02816_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10810__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09008__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06205_ u_cpu.rf_ram.memory\[80\]\[1\] u_cpu.rf_ram.memory\[81\]\[1\] u_cpu.rf_ram.memory\[82\]\[1\]
+ u_cpu.rf_ram.memory\[83\]\[1\] _01706_ _01707_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07019__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07185_ _02758_ _02753_ _02703_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08767__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06136_ _01539_ _01783_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09945__S _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__A2 _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06067_ _01711_ _01714_ _01715_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout401 net406 net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout412 net418 net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07990__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout423 net426 net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout434 net440 net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout445 net447 net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09192__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout456 net458 net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout467 net468 net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09826_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _04544_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07042__I1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06625__S0 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout478 net480 net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout489 net493 net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09757_ _04486_ _04488_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06969_ u_cpu.rf_ram_if.rdata0\[1\] _02599_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11610__CLK net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12736__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10629__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ u_cpu.rf_ram.memory\[140\]\[5\] _03811_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ u_cpu.rf_ram.memory\[122\]\[7\] _04427_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ u_cpu.rf_ram.memory\[15\]\[1\] _03772_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11650_ _00172_ net395 u_cpu.rf_ram.memory\[42\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07213__B _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout30 net32 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout41 net42 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10601_ _05159_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout52 net54 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11581_ _00103_ net214 u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__I0 u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout85 net88 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10532_ _02725_ _05116_ _05118_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xfanout96 net232 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10801__A2 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08823__I _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12116__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10463_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _05072_
+ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12202_ _00716_ net300 u_cpu.rf_ram.memory\[127\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06608__I1 u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10394_ _05034_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10565__A1 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10565__B2 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12133_ _00647_ net61 u_cpu.rf_ram.memory\[134\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07430__A1 u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06233__A2 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09970__A3 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12266__CLK net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07981__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12064_ _00578_ net10 u_cpu.rf_ram.memory\[70\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10317__A1 _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11015_ _05431_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09183__A1 _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06616__S0 _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08930__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12966_ _00092_ net519 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A2 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11917_ _00439_ net220 u_cpu.rf_ram.memory\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07497__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11293__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06544__I0 u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12897_ _01394_ net438 u_cpu.rf_ram.memory\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11424__I _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11848_ _00370_ net102 u_cpu.rf_ram.memory\[66\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09238__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A2 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout235_I net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11779_ _00301_ net273 u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout402_I net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A1 u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06253__I _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12609__CLK net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09410__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__A2 _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _03941_ _03983_ _03991_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ _03210_ _03314_ _03316_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10308__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11633__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09174__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12759__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07872_ _02928_ _03259_ _03265_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07724__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09611_ _04073_ _04389_ _04395_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06823_ _01451_ u_cpu.cpu.bne_or_bge _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06754_ _01634_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout50_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09542_ _04352_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09477__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11783__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07488__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06685_ u_cpu.rf_ram.memory\[108\]\[6\] u_cpu.rf_ram.memory\[109\]\[6\] u_cpu.rf_ram.memory\[110\]\[6\]
+ u_cpu.rf_ram.memory\[111\]\[6\] _02052_ _01506_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _02919_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06160__A1 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09229__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06550__I3 u_cpu.rf_ram.memory\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12139__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08355_ _03563_ _03584_ _03586_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07306_ _02520_ _02526_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08988__A1 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _03493_ _03539_ _03541_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10795__A1 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07237_ _02801_ _02791_ _02790_ _02781_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__12289__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07168_ _02744_ _02738_ _02739_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_106_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07412__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06119_ _01470_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07099_ _02688_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09474__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout220 net221 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11509__I _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout231 net232 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09165__A1 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout242 net243 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout253 net254 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout264 net266 net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout275 net277 net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07715__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout286 net289 net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08912__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09809_ _04511_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout297 net303 net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12820_ _01317_ net100 u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12751_ _01248_ net144 u_cpu.rf_ram.memory\[107\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11702_ _00224_ net387 u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12682_ _01179_ net46 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _00155_ net208 u_cpu.rf_ram.memory\[80\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11027__A2 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08979__A1 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11564_ _05108_ _05777_ _05778_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__A2 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07651__A1 u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _05106_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11495_ _03637_ _05730_ _05737_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10446_ _05064_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11656__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _04800_ _05023_ _05025_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12901__CLK net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07954__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12116_ _00630_ net264 u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05965__A1 _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12047_ _00561_ net17 u_cpu.rf_ram.memory\[73\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08903__A1 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06065__S1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout185_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06390__A1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06780__I3 u_cpu.rf_ram.memory\[123\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout352_I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06517__I0 u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12949_ u_cpu.rf_ram_if.wdata1_r\[1\] net341 u_cpu.rf_ram_if.wdata1_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06470_ u_cpu.rf_ram.memory\[20\]\[4\] u_cpu.rf_ram.memory\[21\]\[4\] u_cpu.rf_ram.memory\[22\]\[4\]
+ u_cpu.rf_ram.memory\[23\]\[4\] _01891_ _02003_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06142__A1 _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11018__A2 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06693__A2 _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08140_ _03418_ _03442_ _03448_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12431__CLK net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__A2 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07237__A4 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ _03341_ _03397_ _03403_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06445__A2 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ u_arbiter.i_wb_cpu_rdt\[1\] _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10529__A1 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08198__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12581__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10434__S _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07945__A2 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06599__I3 u_cpu.rf_ram.memory\[107\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _03052_ _03887_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11329__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07924_ _03301_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10233__I _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07158__B1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09698__A2 _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ u_cpu.rf_ram.memory\[50\]\[6\] _03249_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10701__A1 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08370__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06806_ _01498_ _02438_ _02447_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07786_ _03148_ _03200_ _03208_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__I3 u_cpu.rf_ram.memory\[99\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _04164_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06737_ u_cpu.rf_ram.memory\[16\]\[7\] u_cpu.rf_ram.memory\[17\]\[7\] u_cpu.rf_ram.memory\[18\]\[7\]
+ u_cpu.rf_ram.memory\[19\]\[7\] _02007_ _01518_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11257__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09456_ _04246_ _04297_ _04299_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06668_ _01915_ _02310_ _01663_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06133__B2 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07330__B1 _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09870__A2 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__I3 u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08407_ _03577_ _03610_ _03617_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06684__A2 _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06599_ u_cpu.rf_ram.memory\[104\]\[5\] u_cpu.rf_ram.memory\[105\]\[5\] u_cpu.rf_ram.memory\[106\]\[5\]
+ u_cpu.rf_ram.memory\[107\]\[5\] _02056_ _01624_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09387_ _04246_ _04248_ _04250_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05997__I _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__I _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08338_ _03573_ _03565_ _03574_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10768__A1 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11679__CLK net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08269_ u_cpu.rf_ram.memory\[64\]\[2\] _03530_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ u_cpu.cpu.csr_imm _04949_ _04952_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11280_ _05594_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10231_ u_cpu.cpu.immdec.imm30_25\[2\] _04882_ _04884_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _04892_ _04772_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08189__A2 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07936__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10162_ _04831_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06295__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__A1 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10093_ _04617_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__S1 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11496__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12304__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08361__A2 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06372__A1 _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07452__I _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12803_ _01300_ net415 u_cpu.rf_ram.memory\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10995_ _05419_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08113__A2 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12734_ _01231_ net148 u_cpu.rf_ram.memory\[105\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09861__A2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06675__A2 _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12665_ _01162_ net177 u_cpu.rf_ram.memory\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10208__B1 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11616_ _00138_ net445 u_cpu.rf_ram.memory\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10759__A1 _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12596_ _00021_ net280 u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11420__A2 _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ u_cpu.rf_ram.memory\[23\]\[1\] _05767_ _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11478_ u_cpu.rf_ram.memory\[0\]\[6\] _05722_ _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09377__A1 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ _05055_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11184__A1 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__I _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09129__A1 u_cpu.rf_ram.memory\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ _01618_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10988__I _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07640_ u_cpu.rf_ram.memory\[42\]\[4\] _03110_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07571_ _02946_ _03057_ _03065_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11239__A2 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06522_ _01580_ _02157_ _02166_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09310_ u_cpu.rf_ram.memory\[38\]\[5\] _04197_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10998__A1 _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09852__A2 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06453_ u_cpu.rf_ram.memory\[128\]\[3\] u_cpu.rf_ram.memory\[129\]\[3\] u_cpu.rf_ram.memory\[130\]\[3\]
+ u_cpu.rf_ram.memory\[131\]\[3\] _01747_ _01875_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09241_ _03152_ _03356_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12947__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _04095_ _04104_ _04111_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06384_ _01607_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout13_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08123_ _03422_ _03430_ _03437_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07615__A1 u_cpu.rf_ram.memory\[78\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06418__A2 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11411__A2 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06269__I2 u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08054_ _03347_ _03385_ _03392_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11971__CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07005_ net4 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11175__A1 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06277__S1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10922__A1 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08956_ u_cpu.rf_ram.memory\[136\]\[0\] _03971_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07907_ _03279_ _03294_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11478__A2 _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08887_ _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__A2 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09540__A1 _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07838_ _03228_ _03234_ _03243_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ _03181_ _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ u_cpu.rf_ram.memory\[34\]\[6\] _04325_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10780_ u_cpu.rf_ram.memory\[95\]\[1\] _05284_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09439_ _04283_ _04285_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12450_ _00951_ net482 u_cpu.rf_ram.memory\[113\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05960__S0 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11401_ _05636_ _05671_ _05680_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10138__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07606__A1 u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12381_ _00882_ net472 u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10461__I0 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11332_ _02938_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11263_ u_cpu.rf_ram.memory\[86\]\[3\] _05587_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13002_ _00062_ net525 u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10214_ u_cpu.cpu.immdec.imm30_25\[1\] _04787_ _04682_ _04877_ _04880_ _04881_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08031__A1 u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11194_ _02971_ _05539_ _05544_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10913__A1 u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10145_ u_cpu.rf_ram.memory\[114\]\[7\] _04801_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08582__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09662__I _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10076_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _02709_ _04760_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08334__A2 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08098__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10978_ _05406_ _05401_ _05408_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09834__A2 _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12717_ _01214_ net155 u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07845__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout148_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12648_ _01145_ net144 u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11994__CLK net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout315_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12579_ _01077_ net330 u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11157__A1 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07357__I _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__S1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10904__A1 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ _03875_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _03291_ _04485_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08741_ _03736_ _03832_ _03835_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05953_ u_cpu.rf_ram.memory\[40\]\[0\] u_cpu.rf_ram.memory\[41\]\[0\] u_cpu.rf_ram.memory\[42\]\[0\]
+ u_cpu.rf_ram.memory\[43\]\[0\] _01569_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05884_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08672_ u_cpu.rf_ram.memory\[142\]\[7\] _03782_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07092__I _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06336__B2 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06726__I3 u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07623_ _02879_ _02958_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06887__A2 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07554_ _03054_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06505_ _01646_ _02149_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07485_ u_cpu.rf_ram.memory\[18\]\[4\] _03003_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07836__A1 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06639__A2 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06195__S0 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09224_ u_cpu.rf_ram.memory\[125\]\[1\] _04141_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06436_ _01537_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06436__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09589__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06367_ _02011_ _02012_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09155_ _04099_ _04086_ _04100_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__A2 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08106_ u_cpu.rf_ram.memory\[74\]\[7\] _03409_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08261__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06298_ _01660_ _01944_ _01663_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09086_ _03993_ _04051_ _04053_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08037_ u_cpu.rf_ram.memory\[129\]\[7\] _03371_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11148__A1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__A1 u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09761__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _02707_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10371__A2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _03930_ _03958_ _03961_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06670__S1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09513__A1 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11950_ _00472_ net25 u_cpu.rf_ram.memory\[55\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11320__A1 u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10123__A2 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ u_cpu.rf_ram.memory\[101\]\[6\] _05355_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11881_ _00403_ net185 u_cpu.rf_ram.memory\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10832_ u_cpu.rf_ram.memory\[28\]\[2\] _05318_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10763_ u_cpu.rf_ram.memory\[94\]\[2\] _05275_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__S0 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12502_ _01003_ net490 u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06346__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _05221_ _05199_ _05222_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12433_ _00934_ net233 u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12364_ _00865_ net414 u_cpu.rf_ram.memory\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08252__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11315_ _05619_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12295_ _00796_ net400 u_cpu.rf_ram.memory\[90\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06081__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12642__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ _05562_ _05571_ _05578_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09752__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__A2 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11177_ _05480_ _05526_ _05533_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10362__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10128_ _04160_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_79_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06661__S1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12792__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10059_ _04744_ _04706_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06169__I1 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout265_I net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05916__I1 u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12022__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08736__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10487__B _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout432_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06177__S0 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ _02808_ u_scanchain_local.module_data_in\[63\] _02767_ u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05924__S0 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06221_ _01730_ _01868_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05844__A3 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11378__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06152_ u_cpu.rf_ram.memory\[32\]\[1\] u_cpu.rf_ram.memory\[33\]\[1\] u_cpu.rf_ram.memory\[34\]\[1\]
+ u_cpu.rf_ram.memory\[35\]\[1\] _01590_ _01593_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10050__A1 _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _01517_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10050__B2 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09911_ _02726_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09743__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ _04555_ _04556_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06101__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11550__A1 u_cpu.rf_ram.memory\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10353__A2 _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ u_arbiter.i_wb_cpu_rdt\[1\] _04492_ _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _02608_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08724_ _03631_ _03820_ _03825_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05936_ _01551_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11302__A1 _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06404__S1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08655_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05867_ _01515_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_81_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07606_ u_cpu.rf_ram.memory\[78\]\[0\] _03090_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08586_ u_cpu.rf_ram.memory\[52\]\[1\] _03733_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05798_ u_cpu.cpu.decode.co_ebreak _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07537_ u_cpu.rf_ram.memory\[1\]\[2\] _03043_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12515__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07468_ _02978_ _02988_ _02995_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09207_ u_cpu.rf_ram.memory\[126\]\[2\] _04132_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06419_ _01598_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11369__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07399_ _02876_ u_cpu.rf_ram_if.wdata1_r\[6\] _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09138_ u_cpu.rf_ram.memory\[22\]\[1\] _04086_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08234__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10416__I _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ _04038_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11100_ _05220_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12080_ _00594_ net222 u_cpu.rf_ram.memory\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09734__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08537__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11031_ _05415_ _05433_ _05441_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11541__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06643__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12982_ _00040_ net513 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12045__CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11933_ _00455_ net73 u_cpu.rf_ram.memory\[57\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__B _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _00386_ net105 u_cpu.rf_ram.memory\[64\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10815_ u_cpu.cpu.bufreg.i_sh_signed _04601_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12195__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10100__B _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11795_ _00317_ net18 u_cpu.rf_ram.memory\[74\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06076__I _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _05209_ _05259_ _05265_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07276__A2 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10280__A1 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ u_cpu.rf_ram.memory\[93\]\[3\] _05206_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08225__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12416_ _00917_ net247 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__A1 _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A2 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12347_ _00848_ net452 u_cpu.rf_ram.memory\[118\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06787__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12278_ _00779_ net313 u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09725__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ _05566_ _05553_ _05567_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06539__A1 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11532__A1 u_cpu.rf_ram.memory\[89\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10335__A2 _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout382_I net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06634__S1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _01656_ _02411_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10996__I _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08440_ _03641_ _03625_ _03642_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08700__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08371_ _03167_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] _02871_ u_cpu.cpu.immdec.imm11_7\[0\]
+ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_56_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08464__A1 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12688__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10271__A1 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07253_ _02609_ u_scanchain_local.module_data_in\[60\] _02815_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06570__S0 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09297__I _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06204_ _01704_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07184_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10023__A1 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ u_cpu.rf_ram.memory\[4\]\[1\] u_cpu.rf_ram.memory\[5\]\[1\] u_cpu.rf_ram.memory\[6\]\[1\]
+ u_cpu.rf_ram.memory\[7\]\[1\] _01782_ _01544_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08767__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10574__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06066_ _01555_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout402 net406 net402 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09716__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout413 net418 net413 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout424 net426 net424 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12068__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout435 net439 net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout446 net447 net446 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout457 net458 net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09825_ _04496_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09192__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout468 net469 net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06625__S1 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout479 net483 net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09756_ _02649_ _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06968_ _01471_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08707_ _03746_ _03807_ _03814_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05919_ _01501_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _04176_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ _02536_ _02537_ _02533_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06389__S0 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03621_ _03771_ _03773_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07213__C _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08569_ u_cpu.rf_ram.memory\[53\]\[4\] _03722_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout20 net21 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10600_ _05159_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout42 net96 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08455__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11580_ _00102_ net213 u_cpu.rf_ram.memory\[82\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout75 net76 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10262__A1 u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout86 net88 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_10531_ _05110_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout97 net99 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_109_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10462_ _05073_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12201_ _00715_ net345 u_cpu.rf_ram.memory\[127\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09955__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _03537_ _03231_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10565__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12132_ _00646_ net52 u_cpu.rf_ram.memory\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07430__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09970__A4 _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09707__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12063_ _00577_ net8 u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11514__A1 u_cpu.rf_ram.memory\[100\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11014_ _03182_ _05374_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09183__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06616__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06941__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12965_ _00081_ net522 u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11916_ _00438_ net220 u_cpu.rf_ram.memory\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__A2 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08694__A1 _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12896_ _01393_ net438 u_cpu.rf_ram.memory\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__I _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12830__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _00369_ net100 u_cpu.rf_ram.memory\[66\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11778_ _00300_ net85 u_cpu.rf_ram.memory\[129\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10253__A1 _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout130_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10729_ _04689_ _04631_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout228_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09946__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09845__I _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12210__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07940_ u_cpu.rf_ram.memory\[17\]\[0\] _03315_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11505__A1 u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10308__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07365__I _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07871_ u_cpu.rf_ram.memory\[4\]\[3\] _03263_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07185__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12360__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09610_ u_cpu.rf_ram.memory\[8\]\[3\] _04393_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06232__I0 u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06822_ u_arbiter.i_wb_cpu_dbus_we _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08921__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11928__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ _04352_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06753_ u_cpu.rf_ram.memory\[40\]\[7\] u_cpu.rf_ram.memory\[41\]\[7\] u_cpu.rf_ram.memory\[42\]\[7\]
+ u_cpu.rf_ram.memory\[43\]\[7\] _02027_ _01563_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07488__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09472_ _03103_ _03480_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06684_ _01937_ _02326_ _01596_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08685__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09882__B1 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08423_ _03628_ _03624_ _03629_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ u_cpu.rf_ram.memory\[61\]\[0\] _03585_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07305_ _02856_ _02858_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08285_ u_cpu.rf_ram.memory\[29\]\[0\] _03540_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10795__A2 _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07236_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_30_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06118_ _01763_ _01766_ _01574_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07412__A2 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07098_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_dbus_dat\[28\] _02686_ _02688_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06049_ _01659_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout221 net226 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout232 net512 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09165__A2 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout243 net244 net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout254 net255 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout265 net266 net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout276 net277 net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09808_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _04531_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout287 net289 net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout298 net302 net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06923__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _04433_ _04471_ _04476_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10858__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12750_ _01247_ net144 u_cpu.rf_ram.memory\[107\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11701_ _00223_ net401 u_cpu.rf_ram.memory\[43\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10483__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12681_ _01178_ net46 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06151__A2 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06782__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A1 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11632_ _00154_ net208 u_cpu.rf_ram.memory\[80\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10235__A1 _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ u_cpu.cpu.state.ibus_cyc _05777_ _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11260__I _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06534__S0 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10786__A2 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10514_ _02461_ _02864_ _03270_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_109_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12233__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11494_ u_cpu.rf_ram.memory\[98\]\[4\] _05734_ _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10445_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _05060_
+ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10538__A2 _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__I _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08600__A1 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10376_ u_cpu.rf_ram.memory\[32\]\[0\] _05024_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12115_ _00629_ net264 u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12046_ _00560_ net17 u_cpu.rf_ram.memory\[73\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06914__A1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout178_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__A1 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12948_ _01435_ net334 u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__B1 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12879_ _01376_ net499 u_cpu.rf_ram.memory\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06773__S0 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08419__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout512_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09092__A1 u_cpu.rf_ram.memory\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06525__S0 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08070_ u_cpu.rf_ram.memory\[77\]\[3\] _03401_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07642__A2 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _02641_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09919__A1 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11600__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12726__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10529__A2 _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07309__B _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _03943_ _03971_ _03980_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07095__I _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12876__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ _03215_ _03302_ _03305_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07158__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ _03224_ _03246_ _03253_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10450__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06905__A1 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10701__A2 _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ _02440_ _02442_ _02444_ _02446_ _01613_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ u_cpu.rf_ram.memory\[43\]\[6\] _03203_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12106__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _04339_ _04334_ _04341_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06736_ _01567_ _02377_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06439__I _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08658__A1 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06508__I1 u_cpu.rf_ram.memory\[109\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09455_ u_cpu.rf_ram.memory\[92\]\[0\] _04298_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06667_ u_cpu.rf_ram.memory\[44\]\[6\] u_cpu.rf_ram.memory\[45\]\[6\] u_cpu.rf_ram.memory\[46\]\[6\]
+ u_cpu.rf_ram.memory\[47\]\[6\] _01661_ _02030_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06133__A2 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07330__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06764__S0 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__B2 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08406_ u_cpu.rf_ram.memory\[19\]\[5\] _03613_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09386_ u_cpu.rf_ram.memory\[91\]\[0\] _04249_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12256__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ _01941_ _02241_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08337_ u_cpu.rf_ram.memory\[62\]\[3\] _03571_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10768__A2 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07633__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _03525_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08830__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07219_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _02781_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06692__I0 u_cpu.rf_ram.memory\[120\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08199_ _03413_ _03482_ _03485_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09386__A2 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _04888_ _04894_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06902__I _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11193__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _04828_ _04830_ _04833_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10940__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10092_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _04774_ _04775_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08897__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06777__C _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11255__I _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12802_ _01299_ net415 u_cpu.rf_ram.memory\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08649__A1 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _03086_ _03230_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12733_ _01230_ net120 u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06755__S0 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12664_ _01161_ net197 u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10208__A1 _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11615_ _00137_ net442 u_cpu.rf_ram.memory\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10208__B2 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11623__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12595_ _01093_ net166 u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10759__A2 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11546_ _03620_ _05766_ _05768_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08821__A1 u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06017__C _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11477_ _02978_ _05719_ _05726_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09395__I _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _05054_
+ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09377__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11773__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12899__CLK net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11184__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _04676_ _05010_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10931__A2 _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06060__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout295_I net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12029_ _00543_ net419 u_cpu.rf_ram.memory\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__A1 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout462_I net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07560__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06363__A2 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11165__I _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07570_ u_cpu.rf_ram.memory\[7\]\[6\] _03060_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12279__CLK net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06521_ _02159_ _02161_ _02163_ _02165_ _02072_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07312__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06746__S0 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10998__A2 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _04151_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06452_ _02074_ _02097_ _01743_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09171_ u_cpu.rf_ram.memory\[128\]\[4\] _04108_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06383_ _01599_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08122_ u_cpu.rf_ram.memory\[76\]\[5\] _03433_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07615__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ u_cpu.rf_ram.memory\[139\]\[5\] _03388_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10445__S _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _02463_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07818__I _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07379__A1 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11175__A2 _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08955_ _03969_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07906_ _02616_ _03292_ _03293_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__A1 u_cpu.rf_ram.memory\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ _03052_ _03104_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10686__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ u_cpu.rf_ram.memory\[47\]\[7\] _03232_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09540__A2 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11075__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07768_ _03196_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09507_ _04260_ _04322_ _04329_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06719_ _02342_ _02361_ _01475_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11646__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07303__A1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07699_ _03011_ _03081_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10989__A2 _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09438_ _02482_ _04284_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07854__A2 _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05801__I u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09369_ _04236_ _04237_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__B _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11400_ u_cpu.rf_ram.memory\[27\]\[7\] _05669_ _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05960__S1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12380_ _00881_ net479 u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08803__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11796__CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _05630_ _05620_ _05631_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10610__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _05557_ _05583_ _05588_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13001_ _00061_ net525 u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06417__I0 u_cpu.rf_ram.memory\[120\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10213_ _03278_ _04879_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ u_cpu.rf_ram.memory\[10\]\[2\] _05543_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08031__A2 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06042__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10144_ _04176_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_62_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06432__I3 u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07790__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10075_ _04598_ _04694_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12421__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06079__I _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10977_ u_cpu.rf_ram.memory\[99\]\[2\] _05407_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08098__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09295__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12571__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12716_ _01213_ net155 u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07845__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06499__I3 u_cpu.rf_ram.memory\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12647_ _01144_ net145 u_cpu.rf_ram.memory\[95\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06028__B _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__A2 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12578_ _01076_ net329 u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06656__I0 u_cpu.rf_ram.memory\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11529_ _05753_ _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10452__I1 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout308_I net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08270__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08022__A2 _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06033__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07081__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08740_ u_cpu.rf_ram.memory\[72\]\[1\] _03833_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05952_ _01600_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08469__I _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07373__I _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08671_ _03752_ _03784_ _03792_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11669__CLK net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05883_ _01477_ _01482_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07533__A1 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07622_ _03031_ _03090_ _03099_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12914__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ _03050_ _03053_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06504_ u_cpu.rf_ram.memory\[100\]\[4\] u_cpu.rf_ram.memory\[101\]\[4\] u_cpu.rf_ram.memory\[102\]\[4\]
+ u_cpu.rf_ram.memory\[103\]\[4\] _01934_ _01648_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11093__A1 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ _02974_ _02999_ _03005_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07836__A2 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06195__S1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09223_ _04083_ _04140_ _04142_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06435_ _01852_ _02080_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09154_ u_cpu.rf_ram.memory\[22\]\[6\] _04091_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09589__A2 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06366_ u_cpu.rf_ram.memory\[4\]\[3\] u_cpu.rf_ram.memory\[5\]\[3\] u_cpu.rf_ram.memory\[6\]\[3\]
+ u_cpu.rf_ram.memory\[7\]\[3\] _01782_ _01897_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11396__A2 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08105_ _03352_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09085_ u_cpu.rf_ram.memory\[130\]\[0\] _04052_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06297_ u_cpu.rf_ram.memory\[104\]\[2\] u_cpu.rf_ram.memory\[105\]\[2\] u_cpu.rf_ram.memory\[106\]\[2\]
+ u_cpu.rf_ram.memory\[107\]\[2\] _01661_ _01571_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08261__A2 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__S _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08036_ _03350_ _03373_ _03381_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09210__A1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08013__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__I _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07221__B1 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07072__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12444__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__A2 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10371__A3 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08938_ u_cpu.rf_ram.memory\[49\]\[1\] _03959_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__I _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09513__A2 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _03843_ _03914_ _03916_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__A2 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11320__A2 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12594__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10900_ _05324_ _05352_ _05359_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11880_ _00402_ net181 u_cpu.rf_ram.memory\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ _05311_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _05270_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07827__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12501_ _01002_ net490 u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06186__S1 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ u_cpu.rf_ram.memory\[93\]\[7\] _05197_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12432_ _00933_ net233 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10593__B _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11387__A2 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12363_ _00864_ net414 u_cpu.rf_ram.memory\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08252__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10595__B1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11314_ _05512_ _03328_ _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12294_ _00795_ net400 u_cpu.rf_ram.memory\[90\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11245_ u_cpu.rf_ram.memory\[110\]\[4\] _05575_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07063__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10898__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11176_ u_cpu.rf_ram.memory\[59\]\[4\] _05530_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07763__A1 u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _04805_ _04802_ _04806_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11811__CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07193__I _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09504__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _04708_ _04691_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11311__A2 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05916__I2 u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout160_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11443__I _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout258_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06177__S1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__A1 _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__A1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout425_I net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12317__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05924__S1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06220_ u_cpu.rf_ram.memory\[72\]\[1\] u_cpu.rf_ram.memory\[73\]\[1\] u_cpu.rf_ram.memory\[74\]\[1\]
+ u_cpu.rf_ram.memory\[75\]\[1\] _01867_ _01732_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_106_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05844__A4 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06151_ _01796_ _01798_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09440__A1 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10586__B1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12467__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06272__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06082_ _01540_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09910_ _02706_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06006__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10889__A1 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__B1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ u_arbiter.i_wb_cpu_rdt\[17\] _04546_ _04547_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09743__A2 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11550__A2 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06101__S1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06801__I0 u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ _04499_ _04501_ _04491_ _04502_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07317__B _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06984_ net4 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout73_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ u_cpu.rf_ram.memory\[13\]\[2\] _03824_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05935_ _01583_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11302__A2 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08654_ _03082_ _03370_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05866_ _01514_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07605_ _03088_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _03735_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05797_ u_cpu.cpu.decode.op21 _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11066__A1 _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ _03038_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07467_ u_cpu.rf_ram.memory\[81\]\[5\] _02991_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _04127_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06418_ _01836_ _02063_ _01676_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07398_ _02909_ _02940_ _02941_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11369__A2 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09137_ _03735_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06349_ _01987_ _01989_ _01991_ _01995_ _01768_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08234__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__B1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10041__A2 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09068_ _03998_ _04039_ _04042_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06796__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08019_ _02985_ _03370_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ u_cpu.rf_ram.memory\[105\]\[6\] _05436_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09734__A2 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11984__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12981_ _00039_ net513 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09442__B _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11932_ _00454_ net38 u_cpu.rf_ram.memory\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08170__A1 u_cpu.rf_ram.memory\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11863_ _00385_ net98 u_cpu.rf_ram.memory\[64\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _05221_ _05296_ _05305_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06357__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11794_ _00316_ net165 u_cpu.rf_ram.memory\[77\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__A1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ u_cpu.rf_ram.memory\[97\]\[3\] _05263_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08473__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09668__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10280__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ _05208_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12415_ _00916_ net249 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08225__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10568__B1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12346_ _00847_ net455 u_cpu.rf_ram.memory\[118\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09973__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06787__A2 _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12277_ _00778_ net319 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07036__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11228_ u_cpu.rf_ram.memory\[85\]\[6\] _05558_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09725__A2 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06820__I _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07736__A1 u_cpu.rf_ram.memory\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11532__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11159_ _05482_ _05515_ _05522_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout375_I net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10099__A2 _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08161__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11048__A1 u_cpu.rf_ram.memory\[106\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08370_ _03581_ _03585_ _03594_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ u_cpu.cpu.immdec.imm11_7\[3\] _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_17_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07252_ _02811_ _02813_ _02814_ _02633_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10271__A2 _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08482__I _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06570__S1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06203_ _01698_ _01850_ _01702_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07183_ _02623_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11857__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06134_ _01503_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11220__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06065_ u_cpu.rf_ram.memory\[84\]\[0\] u_cpu.rf_ram.memory\[85\]\[0\] u_cpu.rf_ram.memory\[86\]\[0\]
+ u_cpu.rf_ram.memory\[87\]\[0\] _01712_ _01713_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout403 net405 net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_67_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout414 net415 net414 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout425 net426 net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout436 net439 net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout447 net448 net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09824_ _04542_ _04543_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout458 net459 net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_100_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout469 net470 net469 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09755_ _03282_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06967_ _02587_ _02597_ _02598_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05918_ _01467_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08706_ u_cpu.rf_ram.memory\[140\]\[4\] _03811_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09686_ _04442_ _04429_ _04443_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06898_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] u_cpu.cpu.mem_bytecnt\[1\]
+ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06389__S1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08637_ u_cpu.rf_ram.memory\[15\]\[0\] _03772_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05849_ _01491_ _01492_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11039__A1 u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08568_ _03671_ _03718_ _03724_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout10 net14 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout21 net22 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ u_cpu.rf_ram.memory\[20\]\[6\] _03021_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout32 net41 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout43 net44 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout54 net55 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08499_ _03681_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09652__A1 _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout76 net94 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10530_ _05117_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06561__S1 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10427__I _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _05072_
+ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08207__A2 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12200_ _00714_ net345 u_cpu.rf_ram.memory\[127\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10392_ _04818_ _05024_ _05033_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06608__I3 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12131_ _00645_ net77 u_cpu.rf_ram.memory\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12012__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09707__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12062_ _00576_ net8 u_cpu.rf_ram.memory\[70\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07718__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11514__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11013_ _05417_ _05421_ _05430_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10162__I _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06941__A2 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06792__I2 u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11278__A1 u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12964_ _00070_ net522 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11915_ _00437_ net213 u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12895_ _01392_ net432 u_cpu.rf_ram.memory\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06544__I2 u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06087__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11846_ _00368_ net100 u_cpu.rf_ram.memory\[66\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11777_ _00299_ net84 u_cpu.rf_ram.memory\[129\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09398__I _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10253__A2 _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10728_ _05247_ _05248_ _05252_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10659_ _02905_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout123_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A2 _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12329_ _00830_ net351 u_cpu.rf_ram.memory\[117\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout492_I net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__A1 u_cpu.rf_ram.memory\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ _02921_ _03259_ _03264_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06821_ _02461_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06932__A2 _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09540_ _03327_ _04179_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06752_ _01559_ _02393_ _01533_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10316__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07381__I _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _04264_ _04298_ _04307_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06683_ u_cpu.rf_ram.memory\[96\]\[6\] u_cpu.rf_ram.memory\[97\]\[6\] u_cpu.rf_ram.memory\[98\]\[6\]
+ u_cpu.rf_ram.memory\[99\]\[6\] _01938_ _01593_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10021__B _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09882__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__A2 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09882__B2 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08422_ u_cpu.rf_ram.memory\[5\]\[1\] _03625_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout36_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08353_ _03583_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09634__A1 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07304_ u_cpu.cpu.bufreg.c_r _02857_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11441__A1 _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ _03538_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07235_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ _02740_ _02742_ _02743_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08940__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07948__A1 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06117_ u_cpu.rf_ram.memory\[132\]\[0\] u_cpu.rf_ram.memory\[133\]\[0\] u_cpu.rf_ram.memory\[134\]\[0\]
+ u_cpu.rf_ram.memory\[135\]\[0\] _01764_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07097_ _02687_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ _01693_ _01696_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06460__I _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout200 net201 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout211 net216 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__12185__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout222 net225 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06059__S0 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout233 net235 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout244 net245 net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout255 net256 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_101_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout266 net267 net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09807_ _04496_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout277 net278 net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout288 net289 net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout299 net302 net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07999_ _03357_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09738_ u_cpu.rf_ram.memory\[33\]\[2\] _04475_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08125__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ u_cpu.rf_ram.memory\[122\]\[1\] _04429_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09873__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__B2 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11700_ _00222_ net390 u_cpu.rf_ram.memory\[43\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12680_ _01177_ net46 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11631_ _00153_ net190 u_cpu.rf_ram.memory\[80\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06782__S1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08428__A2 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09625__A1 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11562_ _04600_ _04241_ _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10513_ _04818_ _05096_ _05105_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06534__S1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _03634_ _05730_ _05736_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10444_ _05063_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12528__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10375_ _05022_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08600__A2 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12114_ _00628_ net291 u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06370__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06611__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10106__B _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11499__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12045_ _00559_ net16 u_cpu.rf_ram.memory\[73\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09681__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08364__A1 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06470__S0 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08116__A1 u_cpu.rf_ram.memory\[76\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12947_ u_cpu.rf_ram_if.rtrig0 net285 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09864__A1 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08667__A2 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06517__I2 u_cpu.rf_ram.memory\[114\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__S0 _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__B2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12878_ _01375_ net496 u_cpu.rf_ram.memory\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06773__S1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout240_I net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09616__A1 u_cpu.rf_ram.memory\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08419__A2 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11829_ _00351_ net11 u_cpu.rf_ram.memory\[68\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout338_I net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12058__CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06525__S1 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06150__I0 u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07020_ u_arbiter.i_wb_cpu_rdt\[0\] _02634_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09919__A2 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06453__I1 u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ u_cpu.rf_ram.memory\[136\]\[7\] _03969_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07922_ u_cpu.rf_ram.memory\[16\]\[1\] _03303_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08355__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06205__I1 u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07853_ u_cpu.rf_ram.memory\[50\]\[5\] _03249_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06804_ _01724_ _02445_ _01702_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06461__S0 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__B _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07784_ _03146_ _03200_ _03207_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08107__A1 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06735_ u_cpu.rf_ram.memory\[20\]\[7\] u_cpu.rf_ram.memory\[21\]\[7\] u_cpu.rf_ram.memory\[22\]\[7\]
+ u_cpu.rf_ram.memory\[23\]\[7\] _01570_ _02003_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09523_ u_cpu.rf_ram.memory\[117\]\[2\] _04340_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09855__A1 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08658__A2 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06508__I2 u_cpu.rf_ram.memory\[110\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09454_ _04296_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06669__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06666_ _01634_ _02308_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08935__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06764__S1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08405_ _03575_ _03609_ _03616_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09385_ _04247_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06597_ u_cpu.rf_ram.memory\[108\]\[5\] u_cpu.rf_ram.memory\[109\]\[5\] u_cpu.rf_ram.memory\[110\]\[5\]
+ u_cpu.rf_ram.memory\[111\]\[5\] _02052_ _01827_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08336_ _03340_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06455__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ _03498_ _03526_ _03529_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06141__I0 u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07218_ _02786_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ u_cpu.rf_ram.memory\[67\]\[1\] _03483_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07149_ _02729_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11575__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ _04832_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12820__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10091_ _04773_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10153__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12970__CLK net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__I _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12801_ _01298_ net415 u_cpu.rf_ram.memory\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10993_ _05417_ _05402_ _05418_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08845__I _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12732_ _01229_ net120 u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12200__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06755__S1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12663_ _01160_ net197 u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11614_ _00136_ net441 u_cpu.rf_ram.memory\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06365__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10208__A2 _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05883__A2 _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12594_ _01092_ net174 u_cpu.rf_ram.memory\[109\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09074__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11545_ u_cpu.rf_ram.memory\[23\]\[0\] _05767_ _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08821__A2 _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06832__A1 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11918__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ u_cpu.rf_ram.memory\[0\]\[5\] _05722_ _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10427_ _05047_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _04774_ u_arbiter.i_wb_cpu_rdt\[19\] _04619_ _05009_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10392__A1 _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06060__A2 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _04599_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__I _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12028_ _00542_ net224 u_cpu.rf_ram.memory\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout190_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout288_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06899__A1 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10695__A2 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__A2 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout455_I net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09837__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06520_ _01683_ _02164_ _01687_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08755__I _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07312__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06746__S1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06451_ _01958_ _02087_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06371__I0 u_cpu.rf_ram.memory\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09170_ _04093_ _04104_ _04110_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06382_ u_cpu.rf_ram.memory\[40\]\[3\] u_cpu.rf_ram.memory\[41\]\[3\] u_cpu.rf_ram.memory\[42\]\[3\]
+ u_cpu.rf_ram.memory\[43\]\[3\] _02027_ _01601_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09065__A2 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _03420_ _03429_ _03436_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08812__A2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ _03344_ _03384_ _03391_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07100__S _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07003_ _02610_ _02626_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__S _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12993__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08954_ _03969_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07905_ _03273_ _02619_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08885_ _03729_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08879__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07000__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06434__S0 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10686__A2 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07836_ _03226_ _03234_ _03242_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12223__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07767_ _03051_ _03100_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09506_ u_cpu.rf_ram.memory\[34\]\[5\] _04325_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06718_ _01958_ _02351_ _02360_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_38_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07698_ _03150_ _03135_ _03151_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08500__A1 u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06737__S1 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06649_ u_cpu.rf_ram.memory\[16\]\[6\] u_cpu.rf_ram.memory\[17\]\[6\] u_cpu.rf_ram.memory\[18\]\[6\]
+ u_cpu.rf_ram.memory\[19\]\[6\] _02007_ _01518_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09437_ _02478_ _04282_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06362__I0 u_cpu.rf_ram.memory\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11091__I _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09368_ _04233_ _04232_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09056__A2 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08319_ u_cpu.rf_ram.memory\[63\]\[6\] _03556_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09299_ u_cpu.rf_ram.memory\[38\]\[0\] _04194_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08803__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11330_ u_cpu.rf_ram.memory\[88\]\[4\] _05626_ _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10071__B1 _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06665__I1 u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10610__A2 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11261_ u_cpu.rf_ram.memory\[86\]\[2\] _05587_ _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13000_ _00060_ net526 u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10212_ _04281_ _04878_ _02618_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11192_ _05538_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10143_ _04816_ _04803_ _04817_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06042__A2 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08319__A1 u_cpu.rf_ram.memory\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07744__I _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07790__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10074_ _02522_ _04699_ _04758_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10677__A2 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07542__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09819__A1 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10976_ _05400_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12715_ _01212_ net134 u_cpu.rf_ram.memory\[104\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12646_ _01143_ net146 u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09047__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12866__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12577_ _01075_ net329 u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07919__I _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06656__I1 u_cpu.rf_ram.memory\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ _03627_ _05754_ _05757_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11890__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _05634_ _05707_ _05715_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06033__A2 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07230__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07081__I1 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07781__A2 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05951_ _01551_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10117__A1 _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ u_cpu.rf_ram.memory\[142\]\[6\] _03787_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05882_ u_cpu.rf_ram.memory\[16\]\[0\] u_cpu.rf_ram.memory\[17\]\[0\] u_cpu.rf_ram.memory\[18\]\[0\]
+ u_cpu.rf_ram.memory\[19\]\[0\] _01529_ _01530_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10668__A2 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08730__A1 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07533__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07621_ u_cpu.rf_ram.memory\[78\]\[7\] _03088_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _03052_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08485__I _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05902__I u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06503_ _01499_ _02119_ _02128_ _02147_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07483_ u_cpu.rf_ram.memory\[18\]\[3\] _03003_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11093__A2 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06434_ u_cpu.rf_ram.memory\[80\]\[3\] u_cpu.rf_ram.memory\[81\]\[3\] u_cpu.rf_ram.memory\[82\]\[3\]
+ u_cpu.rf_ram.memory\[83\]\[3\] _01706_ _01965_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ u_cpu.rf_ram.memory\[125\]\[0\] _04141_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09038__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09153_ _03751_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06365_ _01538_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10456__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08104_ _03424_ _03411_ _03425_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06647__I1 u_cpu.rf_ram.memory\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09084_ _04050_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06296_ _01941_ _01942_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08035_ u_cpu.rf_ram.memory\[129\]\[6\] _03376_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13021__CLK net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08549__A1 u_cpu.rf_ram.memory\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10356__A1 _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09210__A2 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07221__A1 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09986_ _03277_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07772__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08937_ _03925_ _03958_ _03960_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06407__S0 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08868_ u_cpu.rf_ram.memory\[138\]\[0\] _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ _03181_ _03231_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08799_ u_cpu.rf_ram.memory\[71\]\[6\] _03868_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _05204_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11763__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10761_ _05202_ _05271_ _05274_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12500_ _01001_ net491 u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10692_ _05220_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12431_ _00932_ net233 u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12119__CLK net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12362_ _00863_ net423 u_cpu.rf_ram.memory\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10595__B2 _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ _02906_ _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06263__A2 _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12293_ _00794_ net380 u_cpu.rf_ram.memory\[90\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12269__CLK net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11244_ _05560_ _05571_ _05577_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10347__A1 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10198__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06015__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07063__I1 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ _05478_ _05526_ _05532_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10898__A2 _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10126_ u_cpu.rf_ram.memory\[114\]\[1\] _04803_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__B _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10057_ _03275_ u_arbiter.i_wb_cpu_rdt\[10\] _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06169__I3 u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05916__I3 u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout153_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10959_ _05322_ _05388_ _05395_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06039__B _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__A2 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__I3 u_cpu.rf_ram.memory\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout320_I net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12629_ _01126_ net205 u_cpu.rf_ram.memory\[97\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout418_I net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__B1 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06150_ u_cpu.rf_ram.memory\[36\]\[1\] u_cpu.rf_ram.memory\[37\]\[1\] u_cpu.rf_ram.memory\[38\]\[1\]
+ u_cpu.rf_ram.memory\[39\]\[1\] _01797_ _01586_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09440__A2 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06081_ _01704_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10008__C _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11636__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__A2 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _04544_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__A2 _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__A1 u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ _02651_ _04489_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06801__I1 u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06983_ _02599_ _02597_ _02607_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ _03819_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05934_ _01514_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout66_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11786__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08703__A1 _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08653_ _03647_ _03772_ _03781_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05865_ u_cpu.raddr\[0\] _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07604_ _03088_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05796_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08584_ _02912_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09104__I _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ _02915_ _03039_ _03042_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11066__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10813__A2 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07466_ _02976_ _02987_ _02994_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09205_ _04088_ _04128_ _04131_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06417_ u_cpu.rf_ram.memory\[120\]\[3\] u_cpu.rf_ram.memory\[121\]\[3\] u_cpu.rf_ram.memory\[122\]\[3\]
+ u_cpu.rf_ram.memory\[123\]\[3\] _01673_ _01837_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ u_cpu.rf_ram.memory\[82\]\[5\] _02922_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09136_ _04083_ _04085_ _04087_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06348_ _01992_ _01994_ _01574_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12411__CLK net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09431__A2 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ u_cpu.rf_ram.memory\[131\]\[1\] _04040_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06279_ _01598_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _03369_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12561__CLK net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08942__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _04605_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12980_ _00038_ net513 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09498__A2 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11931_ _00453_ net70 u_cpu.rf_ram.memory\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09442__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11544__I _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08170__A2 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06181__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11862_ _00384_ net102 u_cpu.rf_ram.memory\[64\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ u_cpu.rf_ram.memory\[96\]\[7\] _05294_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11793_ _00315_ net167 u_cpu.rf_ram.memory\[77\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10804__A2 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10744_ _05205_ _05259_ _05264_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10675_ _02925_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12414_ _00915_ net249 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12091__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10568__A1 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11659__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12345_ _00846_ net350 u_cpu.rf_ram.memory\[118\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12904__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09684__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06787__A3 _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _00777_ net316 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05995__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11227_ _05217_ _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07036__I1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06322__B _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08933__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11158_ u_cpu.rf_ram.memory\[84\]\[5\] _05518_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06041__C _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10109_ _04790_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11089_ u_cpu.rf_ram.memory\[83\]\[3\] _05476_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09489__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11296__A2 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout270_I net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout368_I net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08161__A2 _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout535_I net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09110__A1 u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ u_cpu.cpu.immdec.imm11_7\[4\] _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12434__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _02783_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07672__A1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06202_ u_cpu.rf_ram.memory\[88\]\[1\] u_cpu.rf_ram.memory\[89\]\[1\] u_cpu.rf_ram.memory\[90\]\[1\]
+ u_cpu.rf_ram.memory\[91\]\[1\] _01699_ _01700_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10008__B1 _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _02756_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09413__A2 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ _01773_ _01776_ _01778_ _01780_ _01490_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07424__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06078__I2 u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11220__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12584__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06064_ _01562_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09177__A1 u_cpu.rf_ram.memory\[128\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout404 net405 net404 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout415 net417 net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout426 net427 net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout437 net439 net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09823_ u_arbiter.i_wb_cpu_rdt\[12\] _04533_ _04534_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout448 net449 net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout459 net460 net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10731__A1 _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09754_ _04485_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06966_ _02583_ u_cpu.rf_ram_if.rdata1\[6\] _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08705_ _03743_ _03807_ _03813_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05917_ _01560_ _01565_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09685_ u_cpu.rf_ram.memory\[122\]\[6\] _04434_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06897_ _02505_ _02534_ _02535_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08636_ _03770_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05848_ _01476_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06163__A1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11039__A2 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08567_ u_cpu.rf_ram.memory\[53\]\[3\] _03722_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09101__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout11 net13 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout22 net42 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07518_ _02945_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout33 net36 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout44 net55 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_39_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08498_ _03681_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout55 net95 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09652__A2 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout66 net76 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07663__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout77 net81 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07449_ u_cpu.rf_ram.memory\[21\]\[7\] _02965_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout88 net92 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11801__CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout99 net104 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10460_ _05047_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09119_ _02933_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06218__A2 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07415__A1 u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ u_cpu.rf_ram.memory\[32\]\[7\] _05022_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12130_ _00644_ net259 u_cpu.rf_ram.memory\[135\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11951__CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__C _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__A1 u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09168__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12061_ _00575_ net8 u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09009__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ u_cpu.rf_ram.memory\[79\]\[7\] _05419_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10722__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12307__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__A2 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06796__C _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06792__I3 u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12963_ _00059_ net522 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09340__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08143__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11914_ _00436_ net375 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12894_ _01391_ net432 u_cpu.rf_ram.memory\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06544__I3 u_cpu.rf_ram.memory\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _00367_ net100 u_cpu.rf_ram.memory\[66\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _00298_ net84 u_cpu.rf_ram.memory\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07654__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10727_ _04720_ _05251_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06457__A2 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11450__A2 _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10658_ _04081_ _05185_ _05194_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A2 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__A2 _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09946__A3 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10589_ _05151_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12328_ _00829_ net351 u_cpu.rf_ram.memory\[117\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11449__I _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10961__A1 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09159__A1 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12259_ _00760_ net355 u_cpu.rf_ram.memory\[37\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__A1 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout485_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10713__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _02460_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__I2 u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__I _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06751_ u_cpu.rf_ram.memory\[32\]\[7\] u_cpu.rf_ram.memory\[33\]\[7\] u_cpu.rf_ram.memory\[34\]\[7\]
+ u_cpu.rf_ram.memory\[35\]\[7\] _01745_ _02024_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11269__A2 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10316__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09331__A1 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08134__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ u_cpu.rf_ram.memory\[92\]\[7\] _04296_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06682_ _01656_ _02324_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06145__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10021__C _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09882__A2 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _03627_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08352_ _03583_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05910__I _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout29_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07303_ _02480_ _02850_ _02851_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07645__A1 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10528__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11441__A2 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _03538_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07234_ _02724_ _02798_ _02799_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _02684_ u_scanchain_local.module_data_in\[45\] _02730_ u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06116_ _01721_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08070__A1 u_cpu.rf_ram.memory\[77\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07096_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_dbus_dat\[27\] _02686_ _02687_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__A1 _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06047_ u_cpu.rf_ram.memory\[92\]\[0\] u_cpu.rf_ram.memory\[93\]\[0\] u_cpu.rf_ram.memory\[94\]\[0\]
+ u_cpu.rf_ram.memory\[95\]\[0\] _01694_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06620__A2 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout201 net202 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout212 net215 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout223 net225 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10165__C1 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout234 net235 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout245 net257 net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout256 net257 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09806_ _04529_ _04530_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout267 net278 net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout278 net305 net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout289 net290 net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07998_ _03357_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _04470_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06949_ _02585_ u_cpu.rf_ram.rdata\[1\] _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11094__I _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10212__B _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09322__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08125__A2 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06188__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06136__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09668_ _04157_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09873__A2 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08619_ _03628_ _03758_ _03761_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09599_ _04350_ _04378_ _04387_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _00152_ net187 u_cpu.rf_ram.memory\[80\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05820__I _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11432__A2 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ _03646_ _05767_ _05776_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10438__I _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10512_ u_cpu.rf_ram.memory\[30\]\[7\] _05094_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11492_ u_cpu.rf_ram.memory\[98\]\[3\] _05734_ _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10443_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _05060_
+ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11196__A1 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _05022_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10943__A1 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12113_ _00627_ net291 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06611__A2 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12044_ _00558_ net33 u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08364__A2 _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__I _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06375__A1 _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__B _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__S1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11847__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__A1 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06098__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12946_ _01434_ net320 u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11120__A1 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09864__A2 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__S1 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06678__A2 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12877_ _01374_ net496 u_cpu.rf_ram.memory\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11828_ _00350_ net18 u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout233_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11759_ _00281_ net453 u_cpu.rf_ram.memory\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout400_I net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08052__A1 _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10934__A1 u_cpu.rf_ram.memory\[103\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06453__I2 u_cpu.rf_ram.memory\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08970_ _03941_ _03971_ _03979_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07921_ _03210_ _03302_ _03304_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12622__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08355__A2 _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__I2 u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__I _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07852_ _03222_ _03245_ _03252_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06803_ u_cpu.rf_ram.memory\[76\]\[7\] u_cpu.rf_ram.memory\[77\]\[7\] u_cpu.rf_ram.memory\[78\]\[7\]
+ u_cpu.rf_ram.memory\[79\]\[7\] _01725_ _01726_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07783_ u_cpu.rf_ram.memory\[43\]\[5\] _03203_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07325__C _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06461__S1 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12772__CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09522_ _04333_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06734_ _01719_ _02375_ _02001_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__A1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09855__A2 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ _04296_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06665_ u_cpu.rf_ram.memory\[40\]\[6\] u_cpu.rf_ram.memory\[41\]\[6\] u_cpu.rf_ram.memory\[42\]\[6\]
+ u_cpu.rf_ram.memory\[43\]\[6\] _02027_ _01563_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08404_ u_cpu.rf_ram.memory\[19\]\[4\] _03613_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09384_ _04247_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12002__CLK net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06596_ _01937_ _02239_ _01596_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09112__I _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07618__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08335_ _03570_ _03565_ _03572_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11414__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08291__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08266_ u_cpu.rf_ram.memory\[64\]\[1\] _03527_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07094__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__I1 u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07217_ _02634_ u_scanchain_local.module_data_in\[54\] _02785_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12152__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11178__A1 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03408_ _03482_ _03484_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08043__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ _02628_ _02702_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07079_ _02676_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09782__I _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10090_ _02707_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08346__A2 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09543__A1 u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10153__A2 _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12800_ _01297_ net413 u_cpu.rf_ram.memory\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10992_ u_cpu.rf_ram.memory\[99\]\[7\] _05400_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11102__A1 _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12731_ _01228_ net124 u_cpu.rf_ram.memory\[79\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12662_ _01159_ net197 u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _00135_ net382 u_cpu.rf_ram.memory\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07609__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11405__A2 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12593_ _01091_ net171 u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11544_ _05765_ _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08282__A1 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11475_ _02976_ _05718_ _05725_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06683__I2 u_cpu.rf_ram.memory\[98\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06381__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _05053_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08034__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12645__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10916__A1 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10357_ _02709_ _02648_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09692__I _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10288_ _04947_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08337__A2 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12027_ _00541_ net224 u_cpu.rf_ram.memory\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11341__A1 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout183_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12025__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09837__A2 _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12929_ _01425_ net378 u_cpu.rf_ram.memory\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout350_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07848__A1 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout448_I net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ _02089_ _02091_ _02093_ _02095_ _01982_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_61_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__I1 u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _01568_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08120_ u_cpu.rf_ram.memory\[76\]\[4\] _03433_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08771__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08051_ u_cpu.rf_ram.memory\[139\]\[4\] _03388_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06823__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__I2 u_cpu.rf_ram.memory\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07387__I _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05882__I0 u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07002_ _02613_ _02620_ _02625_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06291__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06224__C _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08576__A2 _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06131__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08953_ _03327_ _03887_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08328__A2 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07904_ _02557_ _03290_ _03291_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ _03861_ _03915_ _03924_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07835_ u_cpu.rf_ram.memory\[47\]\[6\] _03237_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07000__A2 _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06434__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ _03150_ _03186_ _03195_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09505_ _04258_ _04321_ _04328_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07839__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06717_ _02353_ _02355_ _02357_ _02359_ _01982_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_53_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ u_cpu.rf_ram.memory\[45\]\[7\] _03133_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12518__CLK net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07303__A3 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08500__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09436_ _02480_ _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06648_ _01890_ _02290_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06511__A1 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05945__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09367_ u_cpu.cpu.mem_bytecnt\[1\] _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06579_ u_cpu.rf_ram.memory\[44\]\[5\] u_cpu.rf_ram.memory\[45\]\[5\] u_cpu.rf_ram.memory\[46\]\[5\]
+ u_cpu.rf_ram.memory\[47\]\[5\] _01805_ _02030_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11399__A1 _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08318_ _03507_ _03553_ _03560_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08681__I _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09298_ _04192_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10071__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08249_ u_cpu.rf_ram.memory\[65\]\[2\] _03518_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10071__B2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08016__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11260_ _05582_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11692__CLK net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09764__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _02614_ _02615_ _02463_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _02969_ _05539_ _05542_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06417__I2 u_cpu.rf_ram.memory\[122\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06578__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11571__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ u_cpu.rf_ram.memory\[114\]\[6\] _04808_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06042__A3 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09445__C _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08319__A2 _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10073_ _04720_ _04757_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10126__A2 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09819__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06750__A1 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12198__CLK net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10975_ _05204_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12714_ _01211_ net134 u_cpu.rf_ram.memory\[104\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06309__C _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12645_ _01142_ net152 u_cpu.rf_ram.memory\[95\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09687__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12576_ _01074_ net329 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11527_ u_cpu.rf_ram.memory\[89\]\[1\] _05755_ _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08007__A1 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11458_ u_cpu.rf_ram.memory\[24\]\[6\] _05710_ _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10409_ u_cpu.rf_ram.memory\[31\]\[6\] _05039_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11389_ _05669_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11562__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout398_I net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09507__A1 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ _01598_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11314__A1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10117__A2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05881_ _01517_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _03029_ _03090_ _03098_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__A1 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07551_ _02959_ _03051_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10310__B _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _01795_ _02137_ _02146_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ _02971_ _02999_ _03004_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _04139_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06433_ _01698_ _02078_ _01963_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09152_ _04097_ _04086_ _04098_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout11_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06364_ _01999_ _02002_ _02005_ _02009_ _01490_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08103_ u_cpu.rf_ram.memory\[74\]\[6\] _03416_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08797__A2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06295_ u_cpu.rf_ram.memory\[108\]\[2\] u_cpu.rf_ram.memory\[109\]\[2\] u_cpu.rf_ram.memory\[110\]\[2\]
+ u_cpu.rf_ram.memory\[111\]\[2\] _01549_ _01827_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09083_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06647__I2 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06352__S0 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12960__CLK net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06235__B _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08034_ _03347_ _03373_ _03380_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10472__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11553__A1 _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09985_ _02542_ _04601_ _04675_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08936_ u_cpu.rf_ram.memory\[49\]\[0\] _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06407__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08867_ _03913_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06032__I0 u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07818_ _03230_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08676__I _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ _03857_ _03865_ _03872_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11908__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _03184_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ u_cpu.rf_ram.memory\[94\]\[1\] _05272_ _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12490__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09419_ _04253_ _04267_ _04272_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ _02949_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12430_ _00931_ net49 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08237__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08788__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12361_ _00862_ net423 u_cpu.rf_ram.memory\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06343__S0 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10595__A2 _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11312_ _05568_ _05608_ _05617_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12292_ _00793_ net398 u_cpu.rf_ram.memory\[90\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11243_ u_cpu.rf_ram.memory\[110\]\[3\] _05575_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10347__A2 _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11174_ u_cpu.rf_ram.memory\[59\]\[3\] _05530_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _04157_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10181__I _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ _02707_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08712__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06723__A1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10958_ u_cpu.rf_ram.memory\[104\]\[4\] _05392_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__A3 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10889_ _05309_ _05351_ _05353_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06582__S0 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12628_ _01125_ net159 u_cpu.rf_ram.memory\[97\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08228__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10035__A1 _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A1 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__B2 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A2 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout313_I net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12559_ _01057_ net308 u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10586__A2 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06080_ _01724_ _01727_ _01728_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12213__CLK net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__A1 _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08400__A1 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06262__I0 u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _04486_ _04500_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__A2 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06982_ u_cpu.rf_ram_if.rdata0\[7\] _02602_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _03628_ _03820_ _03823_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05933_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ u_cpu.rf_ram.memory\[15\]\[7\] _03770_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05864_ _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06714__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10510__A2 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05913__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ _03083_ _03087_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08583_ _03730_ _03732_ _03734_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05795_ _01442_ _01445_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07534_ u_cpu.rf_ram.memory\[1\]\[1\] _03040_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__A1 u_cpu.rf_ram.memory\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07465_ u_cpu.rf_ram.memory\[81\]\[4\] _02991_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10467__S _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09204_ u_cpu.rf_ram.memory\[126\]\[1\] _04129_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06416_ _01667_ _02061_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07396_ _02939_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ u_cpu.rf_ram.memory\[22\]\[0\] _04086_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09967__A1 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11369__A4 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06347_ u_cpu.rf_ram.memory\[132\]\[2\] u_cpu.rf_ram.memory\[133\]\[2\] u_cpu.rf_ram.memory\[134\]\[2\]
+ u_cpu.rf_ram.memory\[135\]\[2\] _01993_ _01765_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10577__A2 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09066_ _03993_ _04039_ _04041_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06278_ _01629_ _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09719__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ _02892_ _02962_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11526__A1 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10329__A2 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__I _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09195__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11097__I _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09968_ _04602_ _02648_ _04659_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11730__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12856__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ _03930_ _03946_ _03949_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09899_ _04440_ _04586_ _04593_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11930_ _00452_ net72 u_cpu.rf_ram.memory\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06919__I _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06705__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11861_ _00383_ net102 u_cpu.rf_ram.memory\[64\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11880__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10812_ _05218_ _05296_ _05304_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08458__A1 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11792_ _00314_ net167 u_cpu.rf_ram.memory\[77\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10265__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ u_cpu.rf_ram.memory\[97\]\[2\] _05263_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12236__CLK net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10674_ _05205_ _05198_ _05207_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12413_ _00914_ net247 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10568__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12344_ _00845_ net350 u_cpu.rf_ram.memory\[118\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08630__A1 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12275_ _00776_ net314 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11517__A1 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05995__A2 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ _05564_ _05553_ _05565_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__A2 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11157_ _05480_ _05514_ _05521_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06944__A1 _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10740__A2 _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _04622_ _04652_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11088_ _05208_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10879__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10039_ _04708_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout263_I net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__A2 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__A1 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09110__A2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout430_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout528_I net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06555__S0 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ _02703_ _02812_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07672__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06201_ _01693_ _01848_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10008__A1 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10008__B2 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07181_ _02609_ u_scanchain_local.module_data_in\[48\] _02625_ u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _02755_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_30_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12729__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06307__S0 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06132_ _01528_ _01779_ _01534_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07424__A2 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06078__I3 u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06063_ _01502_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07395__I _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11508__A1 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout405 net406 net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07188__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout416 net418 net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout427 net428 net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09822_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _04531_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08924__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout438 net439 net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout449 net450 net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10731__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ _03280_ _04484_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06965_ _02474_ u_cpu.rf_ram.rdata\[6\] _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12109__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08704_ u_cpu.rf_ram.memory\[140\]\[3\] _03811_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05916_ u_cpu.rf_ram.memory\[8\]\[0\] u_cpu.rf_ram.memory\[9\]\[0\] u_cpu.rf_ram.memory\[10\]\[0\]
+ u_cpu.rf_ram.memory\[11\]\[0\] _01561_ _01564_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09684_ _04173_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06896_ _02505_ _02469_ _02470_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06538__I1 u_cpu.rf_ram.memory\[77\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08635_ _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05847_ _01496_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06794__S0 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ _03668_ _03718_ _03723_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12259__CLK net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__A1 _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout12 net13 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07517_ _03027_ _03016_ _03028_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09101__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__B _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout23 net27 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03550_ _03328_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout34 net35 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06546__S0 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout45 net46 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10798__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout56 net60 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_39_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout67 net69 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07448_ _02950_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A1 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout78 net81 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout89 net92 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ _02902_ u_cpu.rf_ram_if.wdata0_r\[3\] _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_108_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _04073_ _04065_ _04074_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10390_ _04816_ _05024_ _05032_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08612__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _04026_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05818__I _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__A2 _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A2 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12060_ _00574_ net22 u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11011_ _05415_ _05421_ _05429_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06926__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10722__A2 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06926__B2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12962_ _00048_ net521 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10486__A1 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09340__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11913_ _00435_ net375 u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12893_ _01390_ net497 u_cpu.rf_ram.memory\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07351__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__A2 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _00366_ net107 u_cpu.rf_ram.memory\[66\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11775_ _00297_ net91 u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07103__A1 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__A2 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06384__I _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10726_ _04664_ _04791_ _04701_ _04702_ _05250_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08851__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07654__A2 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ u_cpu.rf_ram.memory\[2\]\[7\] _05183_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11776__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10588_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _05107_ _05146_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09946__A4 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10410__A1 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12327_ _00828_ net361 u_cpu.rf_ram.memory\[117\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09159__A2 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12258_ _00759_ net355 u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11209_ u_cpu.rf_ram.memory\[85\]\[0\] _05553_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12189_ _00703_ net261 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06917__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout380_I net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06232__I3 u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06750_ _01629_ _02391_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12401__CLK net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ u_cpu.rf_ram.memory\[100\]\[6\] u_cpu.rf_ram.memory\[101\]\[6\] u_cpu.rf_ram.memory\[102\]\[6\]
+ u_cpu.rf_ram.memory\[103\]\[6\] _01934_ _01543_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_92_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06145__A2 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _02913_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08774__I _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07893__A2 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10229__A1 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _03131_ _03168_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09095__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12551__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07302_ _02536_ _02855_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06294__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08282_ _03537_ _03132_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07645__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ _02749_ u_scanchain_local.module_data_in\[57\] _02788_ u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _02696_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06115_ _01541_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08070__A2 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _02664_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06700__S0 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06046_ _01618_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout202 net206 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout213 net215 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout224 net225 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__B1 _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout235 net245 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__C2 _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout246 net247 net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_60_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09805_ u_arbiter.i_wb_cpu_rdt\[7\] _04512_ _04524_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout257 net306 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout268 net272 net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout279 net284 net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07997_ _03053_ _03356_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09736_ _04431_ _04471_ _04474_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06948_ _02474_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09667_ _04425_ _04428_ _04430_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11649__CLK net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06879_ _02517_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06136__A2 _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07333__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ u_cpu.rf_ram.memory\[9\]\[1\] _03759_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09598_ u_cpu.rf_ram.memory\[121\]\[7\] _04376_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06931__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ u_cpu.rf_ram.memory\[54\]\[4\] _03710_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09086__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__S0 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06418__B _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05990__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11560_ u_cpu.rf_ram.memory\[23\]\[7\] _05765_ _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11799__CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__A2 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08833__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _04816_ _05096_ _05104_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ _03630_ _05730_ _05735_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A2 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10442_ _05062_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__A2 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10373_ _03067_ _03130_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10943__A2 _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12112_ _00626_ net291 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06611__A3 _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12043_ _00557_ net33 u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05992__B _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12424__CLK net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__A1 u_cpu.rf_ram.memory\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12945_ _01433_ net279 u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11120__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12574__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06758__S0 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08594__I _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A2 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12876_ _01373_ net500 u_cpu.rf_ram.memory\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09077__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11827_ _00349_ net19 u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11758_ _00280_ net453 u_cpu.rf_ram.memory\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A1 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10709_ _04891_ _04772_ _05235_ _04670_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout226_I net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11689_ _00211_ net456 u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06438__I0 u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10934__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06453__I3 u_cpu.rf_ram.memory\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ u_cpu.rf_ram.memory\[16\]\[0\] _03303_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__A1 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10698__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09552__A2 _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ u_cpu.rf_ram.memory\[50\]\[4\] _03249_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10698__B2 _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06205__I3 u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10313__B _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07563__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06802_ _01705_ _02443_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12917__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07782_ _03144_ _03199_ _03206_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput2 io_in[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _04160_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06733_ u_cpu.rf_ram.memory\[24\]\[7\] u_cpu.rf_ram.memory\[25\]\[7\] u_cpu.rf_ram.memory\[26\]\[7\]
+ u_cpu.rf_ram.memory\[27\]\[7\] _01746_ _01748_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11111__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__S0 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ _04295_ _03153_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06664_ _01559_ _02306_ _01533_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout41_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07866__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05921__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11941__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08403_ _03573_ _03609_ _03615_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09383_ _02899_ _03197_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__A1 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06595_ u_cpu.rf_ram.memory\[96\]\[5\] u_cpu.rf_ram.memory\[97\]\[5\] u_cpu.rf_ram.memory\[98\]\[5\]
+ u_cpu.rf_ram.memory\[99\]\[5\] _01938_ _01824_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08334_ u_cpu.rf_ram.memory\[62\]\[2\] _03571_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08815__A1 u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ _03493_ _03526_ _03528_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08291__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07216_ _02686_ _02782_ _02784_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08196_ u_cpu.rf_ram.memory\[67\]\[0\] _03483_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11178__A2 _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07147_ _02725_ _02727_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06054__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12447__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_dbus_dat\[20\] _02671_ _02676_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ _01598_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12597__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10153__A3 _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06199__I _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09719_ _04433_ _04459_ _04464_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10991_ _05220_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12730_ _01227_ net124 u_cpu.rf_ram.memory\[79\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07857__A2 _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09303__I _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12661_ _01158_ net176 u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10449__I _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09059__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11612_ _00134_ net381 u_cpu.rf_ram.memory\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12592_ _01090_ net174 u_cpu.rf_ram.memory\[109\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07609__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08806__A1 u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10613__A1 u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11543_ _05765_ _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08282__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11474_ u_cpu.rf_ram.memory\[0\]\[4\] _05722_ _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11169__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10425_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _05048_
+ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08034__A2 _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10117__C _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _04765_ _05007_ _04701_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06596__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11814__CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__I _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10287_ _04946_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08589__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__I _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12026_ _00540_ net71 u_cpu.rf_ram.memory\[140\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06348__A2 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11341__A2 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11964__CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout176_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12928_ _01424_ net189 u_cpu.rf_ram.memory\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07848__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12859_ _01356_ net335 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__A2 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06371__I2 u_cpu.rf_ram.memory\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06380_ _01589_ _02025_ _01801_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10604__A1 u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout510_I net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09470__A1 u_cpu.rf_ram.memory\[92\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08273__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07668__I _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03341_ _03384_ _03390_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06284__B2 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__I3 u_cpu.rf_ram.memory\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07001_ _02624_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10308__B _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__I _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07233__B1 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09773__A2 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06131__S1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07784__A1 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06587__A2 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _03943_ _03959_ _03968_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout89_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07903_ _02632_ _02623_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08883_ u_cpu.rf_ram.memory\[138\]\[7\] _03913_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07834_ _03224_ _03234_ _03241_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07765_ u_cpu.rf_ram.memory\[41\]\[7\] _03184_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09289__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11096__A1 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ u_cpu.rf_ram.memory\[34\]\[4\] _04325_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06716_ _01724_ _02358_ _01702_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07696_ _02951_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07839__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09435_ _02492_ _02487_ _02485_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06647_ u_cpu.rf_ram.memory\[20\]\[6\] u_cpu.rf_ram.memory\[21\]\[6\] u_cpu.rf_ram.memory\[22\]\[6\]
+ u_cpu.rf_ram.memory\[23\]\[6\] _01891_ _02003_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06511__A2 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05945__S1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09366_ _04233_ _04232_ _04235_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06578_ _01634_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11399__A2 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08317_ u_cpu.rf_ram.memory\[63\]\[5\] _03556_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09461__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08264__A2 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09297_ _04192_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08248_ _03513_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08179_ _03468_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08016__A2 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09793__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10210_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_rdt\[9\] _04774_ _04877_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11020__A1 _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11190_ u_cpu.rf_ram.memory\[10\]\[1\] _05540_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09764__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07775__A1 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ _04173_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11987__CLK net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10072_ _04753_ _04612_ _04701_ _04756_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_27_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06750__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11087__A1 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10974_ _05404_ _05401_ _05405_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12713_ _01210_ net134 u_cpu.rf_ram.memory\[104\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A2 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12644_ _01141_ net147 u_cpu.rf_ram.memory\[95\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10907__I _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12575_ _01073_ net325 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09452__A1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08255__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11526_ _03620_ _05754_ _05756_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11457_ _05632_ _05707_ _05714_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08007__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12762__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _04814_ _05036_ _05043_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11011__A1 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11388_ _05623_ _05670_ _05673_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07766__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _04897_ _04687_ _04865_ _04988_ _04850_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout293_I net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11314__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12009_ _00523_ net56 u_cpu.rf_ram.memory\[142\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05880_ _01515_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10522__B1 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08191__A1 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout460_I net470 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12142__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ _02887_ _02956_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06501_ _02139_ _02141_ _02143_ _02145_ _01642_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10825__A1 u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07481_ u_cpu.rf_ram.memory\[18\]\[2\] _03003_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10089__I _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _04139_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06432_ u_cpu.rf_ram.memory\[88\]\[3\] u_cpu.rf_ram.memory\[89\]\[3\] u_cpu.rf_ram.memory\[90\]\[3\]
+ u_cpu.rf_ram.memory\[91\]\[3\] _01961_ _01700_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12292__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ u_cpu.rf_ram.memory\[22\]\[5\] _04091_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06363_ _02006_ _02008_ _01534_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08246__A2 _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08102_ _03349_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06516__B _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11250__A1 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ _02890_ _04013_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06294_ _01710_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06647__I3 u_cpu.rf_ram.memory\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__B _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06352__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08033_ u_cpu.rf_ram.memory\[129\]\[5\] _03376_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06009__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11002__A1 u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09746__A2 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A1 u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11553__A2 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10552__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09984_ _04672_ _04620_ _04625_ _04673_ _04674_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_44_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _03957_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11305__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06980__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _03913_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ _03051_ _03081_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ u_cpu.rf_ram.memory\[71\]\[5\] _03868_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11383__I _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06732__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11069__A1 u_cpu.rf_ram.memory\[107\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ _03184_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12635__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10816__A1 _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07679_ _03137_ _03134_ _03138_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ u_cpu.rf_ram.memory\[90\]\[2\] _04271_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10690_ _05218_ _05199_ _05219_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _04168_ _04217_ _04224_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12360_ _00861_ net441 u_cpu.rf_ram.memory\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11241__A1 u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10044__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06638__I3 u_cpu.rf_ram.memory\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11311_ u_cpu.rf_ram.memory\[87\]\[7\] _05606_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06343__S1 _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12291_ _00792_ net398 u_cpu.rf_ram.memory\[90\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12015__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11242_ _05557_ _05571_ _05576_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11173_ _05475_ _05526_ _05531_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07212__A3 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10124_ _04800_ _04802_ _04804_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06810__I3 u_cpu.rf_ram.memory\[135\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06971__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ _04740_ _04688_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A1 u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06723__A2 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10107__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10807__A1 u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10957_ _05320_ _05388_ _05394_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09673__A1 u_cpu.rf_ram.memory\[122\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06487__A1 _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10283__A2 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10888_ u_cpu.rf_ram.memory\[101\]\[0\] _05352_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06582__S1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12627_ _01124_ net205 u_cpu.rf_ram.memory\[97\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09425__A1 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08228__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout139_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11232__A1 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A2 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12558_ _01056_ net250 u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11509_ _05741_ _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout306_I net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12489_ _00990_ net242 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07739__A1 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06262__I1 u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ _02599_ _02595_ _02606_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08720_ u_cpu.rf_ram.memory\[13\]\[1\] _03821_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11299__A1 _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05932_ _01466_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08777__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08164__A1 u_cpu.rf_ram.memory\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _03644_ _03772_ _03780_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05863_ _01511_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09900__A2 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07911__A1 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07602_ _03086_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08582_ u_cpu.rf_ram.memory\[52\]\[0\] _03733_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05794_ _01443_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07533_ _02908_ _03039_ _03041_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11471__A1 _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ _02974_ _02987_ _02993_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10274__A2 _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09401__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06573__S1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06415_ u_cpu.rf_ram.memory\[124\]\[3\] u_cpu.rf_ram.memory\[125\]\[3\] u_cpu.rf_ram.memory\[126\]\[3\]
+ u_cpu.rf_ram.memory\[127\]\[3\] _01947_ _01669_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09203_ _04083_ _04128_ _04130_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07395_ _02938_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09416__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09134_ _04084_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12038__CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11223__A1 _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06346_ _01541_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A1 _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ u_cpu.rf_ram.memory\[131\]\[0\] _04040_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06277_ u_cpu.rf_ram.memory\[52\]\[2\] u_cpu.rf_ram.memory\[53\]\[2\] u_cpu.rf_ram.memory\[54\]\[2\]
+ u_cpu.rf_ram.memory\[55\]\[2\] _01630_ _01631_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ _03353_ _03359_ _03368_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12188__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10734__B1 _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _04605_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06953__A2 u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08918_ u_cpu.rf_ram.memory\[137\]\[1\] _03947_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09898_ u_cpu.rf_ram.memory\[113\]\[5\] _04589_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08849_ _03621_ _03902_ _03904_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06705__A2 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07902__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11860_ _00382_ net108 u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ u_cpu.rf_ram.memory\[96\]\[6\] _05299_ _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11791_ _00313_ net167 u_cpu.rf_ram.memory\[77\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06013__S0 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11462__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10742_ _05258_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06935__I u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ u_cpu.rf_ram.memory\[93\]\[2\] _05206_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12412_ _00913_ net465 u_cpu.rf_ram.memory\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07969__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12343_ _00844_ net346 u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12274_ _00775_ net314 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11225_ u_cpu.rf_ram.memory\[85\]\[5\] _05558_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05995__A3 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09981__I _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ u_cpu.rf_ram.memory\[84\]\[4\] _05518_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _02708_ _04789_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11087_ _05475_ _05470_ _05477_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__I _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08146__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10038_ _04625_ _04673_ _04681_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08697__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12950__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06172__A3 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09646__A1 u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout256_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08449__A2 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11989_ _00511_ net419 u_cpu.rf_ram.memory\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06004__S0 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11453__A1 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06555__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout423_I net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ u_cpu.rf_ram.memory\[92\]\[1\] u_cpu.rf_ram.memory\[93\]\[1\] u_cpu.rf_ram.memory\[94\]\[1\]
+ u_cpu.rf_ram.memory\[95\]\[1\] _01694_ _01847_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10008__A2 _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _02753_ _02754_ _02713_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06880__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06307__S1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ u_cpu.rf_ram.memory\[16\]\[1\] u_cpu.rf_ram.memory\[17\]\[1\] u_cpu.rf_ram.memory\[18\]\[1\]
+ u_cpu.rf_ram.memory\[19\]\[1\] _01529_ _01530_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08621__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06062_ _01710_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09891__I _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08385__A1 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout406 net407 net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout417 net418 net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12480__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09821_ _04540_ _04541_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout428 net450 net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout439 net440 net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10830__I _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ _02460_ _04482_ _04483_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout71_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06964_ _02584_ _02595_ _02596_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08703_ _03739_ _03807_ _03812_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05915_ _01563_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09683_ _04440_ _04429_ _04441_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06895_ u_cpu.cpu.immdec.imm31 _02471_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__A2 _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06538__I2 u_cpu.rf_ram.memory\[78\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06699__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05846_ _01471_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06794__S1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10478__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ u_cpu.rf_ram.memory\[53\]\[2\] _03722_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07516_ u_cpu.rf_ram.memory\[20\]\[5\] _03021_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10247__A2 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout13 net14 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_39_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout24 net26 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_08496_ _03679_ _03664_ _03680_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout35 net36 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09131__I _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06546__S1 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout46 net55 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07447_ _02980_ _02967_ _02981_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout57 net60 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout68 net69 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout79 net80 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06871__B2 _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ _02903_ u_cpu.rf_ram_if.wdata1_r\[3\] _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ u_cpu.rf_ram.memory\[12\]\[3\] _04071_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ _01862_ _01975_ _01865_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08612__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11578__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09048_ _03998_ _04027_ _04030_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12823__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ u_cpu.rf_ram.memory\[79\]\[6\] _05424_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08376__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10722__A3 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12973__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05834__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12961_ _00037_ net529 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09876__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08679__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09876__B2 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09750__B u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__S0 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11912_ _00434_ net276 u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10486__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12892_ _01389_ net505 u_cpu.rf_ram.memory\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12203__CLK net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07351__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11843_ _00365_ net107 u_cpu.rf_ram.memory\[66\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__A1 _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11774_ _00296_ net91 u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A1 u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10725_ _05237_ _05249_ _04908_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12353__CLK net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06162__I0 u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08851__A2 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06862__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _04079_ _05185_ _05193_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ _05150_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08603__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07496__I _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12326_ _00827_ net351 u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12257_ _00758_ net360 u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11208_ _05551_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12188_ _00702_ net260 u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10174__A1 _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06917__A2 _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10713__A3 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11139_ u_cpu.rf_ram.memory\[69\]\[6\] _05505_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05976__I0 u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08119__A1 _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout373_I net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06680_ _01692_ _02294_ _02303_ _02322_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_23_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09619__A1 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07180__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ _03581_ _03566_ _03582_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11426__A1 _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09095__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07301_ _02548_ _02854_ _02557_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08281_ _02963_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09886__I _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _02793_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08790__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07163_ _02738_ _02739_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05919__I _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ _01558_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06605__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10401__A2 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07094_ _02683_ _02643_ _02685_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06700__S1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06045_ _01540_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12996__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout203 net204 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10165__A1 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout225 net226 net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10165__B2 _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout236 net245 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout247 net251 net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09804_ u_arbiter.i_wb_cpu_dbus_dat\[7\] _04526_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout258 net262 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout269 net272 net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07996_ _03355_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07581__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ u_cpu.rf_ram.memory\[33\]\[1\] _04472_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06947_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06216__S0 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09666_ u_cpu.rf_ram.memory\[122\]\[0\] _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06878_ _01444_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07333__A2 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08530__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08617_ _03621_ _03758_ _03760_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05829_ _01448_ _01442_ _01460_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _04348_ _04378_ _04386_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06931__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11417__A1 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08548_ _03671_ _03706_ _03712_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09086__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__S1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _03662_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10510_ u_cpu.rf_ram.memory\[30\]\[6\] _05099_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11490_ u_cpu.rf_ram.memory\[98\]\[2\] _05734_ _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _05060_
+ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__B1 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10372_ _05019_ _05020_ _05021_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12111_ _00625_ net282 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13001__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12042_ _00556_ net33 u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__A1 _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12944_ _01432_ net281 u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08521__A1 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06758__S1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12875_ _01372_ net500 u_cpu.rf_ram.memory\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06609__B _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11408__A1 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _00348_ net199 u_cpu.rf_ram.memory\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05886__A2 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09077__A2 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12869__CLK net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11743__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11757_ _00279_ net452 u_cpu.rf_ram.memory\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10631__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10708_ _03084_ _05233_ _05234_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11688_ _00210_ net456 u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06150__I3 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout121_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10639_ _02891_ _03037_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout219_I net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__I _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12309_ _00810_ net487 u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06694__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12249__CLK net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout490_I net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09001__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10380__I _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06446__S0 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07850_ _03220_ _03245_ _03251_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__A2 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ u_cpu.rf_ram.memory\[72\]\[7\] u_cpu.rf_ram.memory\[73\]\[7\] u_cpu.rf_ram.memory\[74\]\[7\]
+ u_cpu.rf_ram.memory\[75\]\[7\] _01694_ _01695_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07781_ u_cpu.rf_ram.memory\[43\]\[4\] _03203_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput3 io_in[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09520_ _04337_ _04334_ _04338_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06732_ _01523_ _02373_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08785__I _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08512__A1 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06749__S1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ _02898_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06663_ u_cpu.rf_ram.memory\[32\]\[6\] u_cpu.rf_ram.memory\[33\]\[6\] u_cpu.rf_ram.memory\[34\]\[6\]
+ u_cpu.rf_ram.memory\[35\]\[6\] _01745_ _02024_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08402_ u_cpu.rf_ram.memory\[19\]\[3\] _03613_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06594_ _01656_ _02237_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09382_ _04151_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout34_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__A2 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08333_ _03564_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08815__A2 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08264_ u_cpu.rf_ram.memory\[64\]\[0\] _03527_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10622__A2 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06141__I3 u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10555__I _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07215_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13024__CLK net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08195_ _03481_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08579__A1 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _02726_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10386__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06054__A2 _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__S0 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07077_ _02675_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ _01672_ _01675_ _01676_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11616__CLK net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10689__A2 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__A1 u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10153__A4 _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ _02932_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09718_ u_cpu.rf_ram.memory\[116\]\[2\] _04463_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08695__I _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _05415_ _05402_ _05416_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08503__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11766__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ u_cpu.rf_ram.memory\[112\]\[2\] _04418_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10310__A1 _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12660_ _01157_ net176 u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09059__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _00133_ net374 u_cpu.rf_ram.memory\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12591_ _01089_ net174 u_cpu.rf_ram.memory\[109\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08806__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11542_ _02963_ _03053_ _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07490__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__A2 _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ _02974_ _05718_ _05724_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10424_ _05052_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10377__A1 _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09231__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__S0 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10355_ _04703_ _04974_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07793__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _02461_ _04945_ _04680_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12025_ _00539_ net61 u_cpu.rf_ram.memory\[140\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07545__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12927_ _01423_ net189 u_cpu.rf_ram.memory\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10301__B2 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout169_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12858_ _01355_ net317 u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11809_ _00331_ net127 u_cpu.rf_ram.memory\[76\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout336_I net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12789_ _01286_ net70 u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06853__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout503_I net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10375__I _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06284__A2 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07000_ net4 _02623_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12071__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11639__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07233__A1 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06667__S0 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07684__I _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07784__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08981__A1 u_cpu.rf_ram.memory\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08951_ u_cpu.rf_ram.memory\[49\]\[7\] _03957_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05795__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07902_ _02495_ _02522_ _03289_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08882_ _03859_ _03915_ _03923_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11789__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ u_cpu.rf_ram.memory\[47\]\[5\] _03237_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ _03148_ _03186_ _03194_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09289__A2 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09404__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05932__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09503_ _04256_ _04321_ _04327_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06715_ u_cpu.rf_ram.memory\[76\]\[6\] u_cpu.rf_ram.memory\[77\]\[6\] u_cpu.rf_ram.memory\[78\]\[6\]
+ u_cpu.rf_ram.memory\[79\]\[6\] _01979_ _01726_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07695_ _03148_ _03135_ _03149_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _02558_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06646_ _01719_ _02288_ _02001_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06362__I3 u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09365_ _04233_ _04232_ _04234_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06577_ u_cpu.rf_ram.memory\[40\]\[5\] u_cpu.rf_ram.memory\[41\]\[5\] u_cpu.rf_ram.memory\[42\]\[5\]
+ u_cpu.rf_ram.memory\[43\]\[5\] _02027_ _01563_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_16_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07859__I _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08316_ _03505_ _03552_ _03559_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12414__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09296_ _03181_ _03453_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07472__A1 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _03498_ _03514_ _03517_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10359__A1 _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _03413_ _03469_ _03472_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09213__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06658__S0 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11020__A2 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _02712_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12564__CLK net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06712__B _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ _04814_ _04803_ _04815_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07775__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08972__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _04748_ _04749_ _04642_ _04661_ _04755_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__A1 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07527__A2 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06003__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11087__A2 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10973_ u_cpu.rf_ram.memory\[99\]\[1\] _05402_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12712_ _01209_ net151 u_cpu.rf_ram.memory\[104\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06502__A3 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12643_ _01140_ net147 u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__B1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12094__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12574_ _01072_ net325 u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09452__A2 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A1 u_cpu.rf_ram.memory\[81\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11525_ u_cpu.rf_ram.memory\[89\]\[0\] _05755_ _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10195__I _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12907__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11456_ u_cpu.rf_ram.memory\[24\]\[5\] _05710_ _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09204__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10407_ u_cpu.rf_ram.memory\[31\]\[5\] _05039_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11387_ u_cpu.rf_ram.memory\[27\]\[1\] _05671_ _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08963__A1 u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10338_ _04989_ _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11931__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10770__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10269_ _04831_ _04822_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12008_ _00522_ net58 u_cpu.rf_ram.memory\[142\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10522__A1 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout286_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08191__A2 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout453_I net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06500_ _01926_ _02144_ _01929_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07480_ _02998_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _01693_ _02076_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06362_ u_cpu.rf_ram.memory\[16\]\[3\] u_cpu.rf_ram.memory\[17\]\[3\] u_cpu.rf_ram.memory\[18\]\[3\]
+ u_cpu.rf_ram.memory\[19\]\[3\] _02007_ _01530_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ _03748_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03422_ _03411_ _03423_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06293_ _01937_ _01939_ _01654_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12587__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ _04011_ _04040_ _04049_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08032_ _03344_ _03372_ _03379_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10061__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09983_ _04598_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10761__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ _03957_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08865_ _03101_ _03887_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06568__I0 u_cpu.rf_ram.memory\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__A1 _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08182__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07816_ _03228_ _03213_ _03229_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06812__S0 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ _03855_ _03864_ _03871_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07747_ _03181_ _03183_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07678_ u_cpu.rf_ram.memory\[45\]\[1\] _03135_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09682__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09417_ _04266_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06496__A2 _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06629_ _02266_ _02268_ _02270_ _02272_ _01982_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_90_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11804__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10029__B1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ u_cpu.rf_ram.memory\[36\]\[4\] _04221_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06248__A2 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ u_cpu.rf_ram.memory\[123\]\[0\] _04182_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11310_ _05566_ _05608_ _05616_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12290_ _00791_ net398 u_cpu.rf_ram.memory\[90\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11954__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09198__A1 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ u_cpu.rf_ram.memory\[110\]\[2\] _05575_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__A1 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08213__I _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ u_cpu.rf_ram.memory\[59\]\[2\] _05530_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10752__A1 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06161__C _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ u_cpu.rf_ram.memory\[114\]\[0\] _04803_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ _04739_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09370__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06803__S0 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09044__I _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10107__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__A2 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10956_ u_cpu.rf_ram.memory\[104\]\[3\] _05392_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09673__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06487__A2 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11480__A2 _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10887_ _05350_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06731__I0 u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12626_ _01123_ net195 u_cpu.rf_ram.memory\[97\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09425__A2 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11232__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12557_ _01055_ net250 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11508_ _03627_ _05742_ _05745_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12488_ _00989_ net242 u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout201_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11439_ _05634_ _05695_ _05703_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06980_ u_cpu.rf_ram_if.rdata0\[6\] _02602_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05931_ _01493_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11299__A2 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11484__I _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__A1 _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08650_ u_cpu.rf_ram.memory\[15\]\[6\] _03775_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05862_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07601_ _03084_ _02892_ _02896_ _03085_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_93_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _03731_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05793_ u_cpu.cpu.branch_op _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07532_ u_cpu.rf_ram.memory\[1\]\[0\] _03040_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A2 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07463_ u_cpu.rf_ram.memory\[81\]\[3\] _02991_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11471__A2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10274__A3 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ u_cpu.rf_ram.memory\[126\]\[0\] _04129_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06414_ _02049_ _02051_ _02054_ _02059_ _01832_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07394_ _02937_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09416__A2 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07427__A1 u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ _04084_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11223__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06345_ _01558_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09064_ _04038_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06276_ _01622_ _01922_ _01626_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08015_ u_cpu.rf_ram.memory\[119\]\[7\] _03357_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06650__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10734__A1 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09966_ _04656_ _04657_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12602__CLK net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _03925_ _03946_ _03948_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09897_ _04438_ _04585_ _04592_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09352__A1 u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ u_cpu.rf_ram.memory\[14\]\[0\] _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__A2 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08779_ _03859_ _03846_ _03860_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10810_ _05215_ _05296_ _05303_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12752__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11790_ _00312_ net167 u_cpu.rf_ram.memory\[77\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09655__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10741_ _05202_ _05259_ _05262_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06469__A2 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__S1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11462__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__I0 u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10672_ _05197_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12411_ _00912_ net485 u_cpu.rf_ram.memory\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07418__A1 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12342_ _00843_ net346 u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10973__A1 u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12132__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12273_ _00774_ net316 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06641__A2 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11224_ _05214_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09591__A1 _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11155_ _05478_ _05514_ _05520_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12282__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10106_ _01448_ _04677_ _04788_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ u_cpu.rf_ram.memory\[83\]\[2\] _05476_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08146__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ _04648_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__A1 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09894__A2 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11988_ _00510_ net223 u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06004__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11453__A2 _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout151_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10939_ _05322_ _05376_ _05383_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout249_I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10110__C1 _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06180__I1 u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12609_ _01106_ net447 u_cpu.rf_ram.memory\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06880__A2 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout416_I net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ _01523_ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07957__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06061_ _01466_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08909__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12625__CLK net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10716__A1 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout407 net408 net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09820_ u_arbiter.i_wb_cpu_rdt\[11\] _04533_ _04534_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08385__A2 _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout418 net428 net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout429 net430 net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_119_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _04236_ _02611_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06963_ _02583_ u_cpu.rf_ram_if.rdata1\[5\] _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08702_ u_cpu.rf_ram.memory\[140\]\[2\] _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08137__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05914_ _01562_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09682_ u_cpu.rf_ram.memory\[122\]\[5\] _04434_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06894_ _02517_ _02532_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _03050_ _03231_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06699__A2 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05845_ _01469_ _01495_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07896__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12005__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08564_ _03717_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09637__A2 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05940__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07515_ _02939_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07648__A1 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout14 net21 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08495_ u_cpu.rf_ram.memory\[57\]\[7\] _03662_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout25 net26 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout36 net40 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout47 net51 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07446_ u_cpu.rf_ram.memory\[21\]\[6\] _02972_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06320__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_91_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12155__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07377_ _02901_ _02921_ _02923_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _02927_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08073__A1 _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06328_ u_cpu.rf_ram.memory\[68\]\[2\] u_cpu.rf_ram.memory\[69\]\[2\] u_cpu.rf_ram.memory\[70\]\[2\]
+ u_cpu.rf_ram.memory\[71\]\[2\] _01725_ _01863_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10955__A1 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11389__I _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ u_cpu.rf_ram.memory\[132\]\[1\] _04028_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06259_ u_cpu.rf_ram.memory\[12\]\[2\] u_cpu.rf_ram.memory\[13\]\[2\] u_cpu.rf_ram.memory\[14\]\[2\]
+ u_cpu.rf_ram.memory\[15\]\[2\] _01570_ _01572_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10707__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09573__A1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08376__A2 _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11380__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _04638_ _04640_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_24_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09325__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12960_ _00026_ net529 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11132__A1 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__A2 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11911_ _00433_ net276 u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06234__S1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12891_ _01388_ net505 u_cpu.rf_ram.memory\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09750__C u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11842_ _00364_ net106 u_cpu.rf_ram.memory\[67\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05850__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07639__A1 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__A2 _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11773_ _00295_ net84 u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ _04623_ _04749_ _04850_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10655_ u_cpu.rf_ram.memory\[2\]\[6\] _05188_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08064__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12648__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10586_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _05144_ _05146_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__A1 _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12325_ _00826_ net454 u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12256_ _00757_ net349 u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11207_ _05551_ _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09564__A1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08367__A2 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12798__CLK net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12187_ _00701_ net260 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11371__A1 _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11138_ _05482_ _05502_ _05509_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout199_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__A1 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08119__A2 _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ u_cpu.rf_ram.memory\[107\]\[5\] _05461_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11123__A1 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A1 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout366_I net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12959__CLKN net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09619__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11426__A2 _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout533_I net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07300_ _02853_ _02543_ _02615_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _03511_ _03527_ _03536_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06302__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07231_ _02797_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07687__I _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07162_ _02738_ _02739_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08055__A1 u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10937__A1 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10327__B _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ _01758_ _01761_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07093_ u_arbiter.i_wb_cpu_rdt\[29\] _02684_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06605__A2 _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06044_ _01581_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09555__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout204 net206 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout215 net216 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout226 net227 net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10165__A2 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11362__A1 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05935__I _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09407__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _04527_ _04528_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout237 net239 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout248 net251 net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07995_ _03084_ _02897_ _03085_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout259 net262 net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_45_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09307__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _04425_ _04471_ _04473_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06946_ u_cpu.rf_ram_if.rtrig1 _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11114__A1 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09858__A2 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09665_ _04427_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06216__S1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06877_ _02512_ _02516_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ u_cpu.rf_ram.memory\[9\]\[0\] _03759_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05828_ u_cpu.cpu.decode.op26 _01449_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06541__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09596_ u_cpu.rf_ram.memory\[121\]\[6\] _04381_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11417__A2 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06931__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10288__I _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08547_ u_cpu.rf_ram.memory\[54\]\[3\] _03710_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ _03336_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07429_ _02913_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _05061_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__B _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09794__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09794__B2 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _05020_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06152__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12110_ _00624_ net293 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09546__A1 _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__A2 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12041_ _00555_ net26 u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09761__B _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09849__A2 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12943_ u_cpu.rf_ram_if.wtrig0 net285 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12874_ _01371_ net502 u_cpu.rf_ram.memory\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11825_ _00347_ net204 u_cpu.rf_ram.memory\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11408__A2 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09987__I _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08891__I _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08285__A1 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11756_ _00278_ net393 u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10707_ u_cpu.cpu.immdec.imm11_7\[1\] _05233_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11687_ _00209_ net464 u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06391__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10638_ _04081_ _05173_ _05182_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09785__A1 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout114_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10862__S _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _05140_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06143__S0 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12308_ _00809_ net197 u_cpu.rf_ram.memory\[92\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06694__S1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12239_ _00014_ net279 u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08131__I _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout483_I net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06446__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06800_ _01711_ _02441_ _01715_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08760__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07780_ _03142_ _03199_ _03205_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07970__I _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 io_in[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_65_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06731_ u_cpu.rf_ram.memory\[28\]\[7\] u_cpu.rf_ram.memory\[29\]\[7\] u_cpu.rf_ram.memory\[30\]\[7\]
+ u_cpu.rf_ram.memory\[31\]\[7\] _01524_ _01525_ _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_92_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09450_ _03272_ _04229_ _04294_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06662_ _01629_ _02304_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ _03570_ _03609_ _03614_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _04245_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06593_ u_cpu.rf_ram.memory\[100\]\[5\] u_cpu.rf_ram.memory\[101\]\[5\] u_cpu.rf_ram.memory\[102\]\[5\]
+ u_cpu.rf_ram.memory\[103\]\[5\] _01934_ _01543_ _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10458__I0 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08332_ _03336_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08276__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout27_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10083__A1 _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08263_ _03525_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06382__S0 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07214_ _02623_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08028__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _03481_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09776__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08579__A2 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07145_ u_cpu.cpu.genblk1.align.ctrl_misal _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_dbus_dat\[19\] _02671_ _02675_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07251__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__S1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06027_ _01610_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__I _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07003__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07978_ _03341_ _03330_ _03342_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09717_ _04458_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06929_ u_cpu.cpu.mem_if.signbit _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08503__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09648_ _04413_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06514__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12493__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09579_ _04350_ _04366_ _04375_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _00132_ net381 u_cpu.rf_ram.memory\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08267__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12590_ _01088_ net174 u_cpu.rf_ram.memory\[109\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__A1 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11541_ _03646_ _05755_ _05764_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06817__A2 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06373__S0 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__A1 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ u_cpu.rf_ram.memory\[0\]\[3\] _05722_ _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08216__I _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07490__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10423_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _05048_
+ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _04970_ _05004_ _05005_ _05006_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06676__S1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09519__A1 u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07276__B _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _02614_ _02542_ _02471_ _02532_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_12024_ _00538_ net63 u_cpu.rf_ram.memory\[140\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11710__CLK net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12926_ _00025_ net292 u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12857_ _01354_ net334 u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12986__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08258__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11808_ _00330_ net127 u_cpu.rf_ram.memory\[76\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12788_ _01285_ net70 u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11739_ _00261_ net433 u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout231_I net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout329_I net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10860__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12216__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07481__A2 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05882__I3 u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06667__S1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12366__CLK net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08981__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _03941_ _03959_ _03967_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__A1 u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05795__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ _03286_ _03288_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08881_ u_cpu.rf_ram.memory\[138\]\[6\] _03918_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07832_ _03222_ _03233_ _03240_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09930__A1 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07763_ u_cpu.rf_ram.memory\[41\]\[6\] _03189_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09502_ u_cpu.rf_ram.memory\[34\]\[3\] _04325_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06714_ _01705_ _02356_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08497__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ u_cpu.rf_ram.memory\[45\]\[6\] _03140_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06249__C _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09433_ u_cpu.cpu.ctrl.i_jump _04242_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06645_ u_cpu.rf_ram.memory\[24\]\[6\] u_cpu.rf_ram.memory\[25\]\[6\] u_cpu.rf_ram.memory\[26\]\[6\]
+ u_cpu.rf_ram.memory\[27\]\[6\] _01746_ _01748_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ _02621_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06576_ _01559_ _02219_ _01801_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10056__A1 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ u_cpu.rf_ram.memory\[63\]\[4\] _03556_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09295_ _04177_ _04182_ _04191_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08246_ u_cpu.rf_ram.memory\[65\]\[1\] _03515_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10851__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09749__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12709__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08177_ u_cpu.rf_ram.memory\[68\]\[1\] _03470_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07128_ _02701_ u_scanchain_local.module_data_in\[39\] _02704_ _02711_ _02625_ u_arbiter.i_wb_cpu_dbus_adr\[2\]
+ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06658__S1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07059_ u_arbiter.i_wb_cpu_rdt\[14\] u_arbiter.i_wb_cpu_dbus_dat\[11\] _02665_ _02666_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08972__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11308__A1 _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06983__A1 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11733__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10070_ _04702_ _04754_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08724__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ _05201_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12711_ _01208_ net151 u_cpu.rf_ram.memory\[104\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10295__B2 _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12642_ _01139_ net148 u_cpu.rf_ram.memory\[95\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12239__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07051__S _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__A1 _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09988__A1 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__B2 _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12573_ _01071_ net325 u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11524_ _05753_ _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A2 _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08660__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11455_ _05630_ _05706_ _05713_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10406_ _04812_ _05035_ _05042_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07215__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _05618_ _05670_ _05672_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06649__S1 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10337_ _04850_ _04990_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08963__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11100__I _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10770__A2 _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10268_ _04923_ _04924_ _04929_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06026__I0 u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12007_ _00521_ net56 u_cpu.rf_ram.memory\[142\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _04862_ _04714_ _04865_ _04866_ _04791_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06577__I1 u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10522__A2 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout181_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06069__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10286__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12909_ _01406_ net196 u_cpu.rf_ram.memory\[98\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout446_I net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ u_cpu.rf_ram.memory\[92\]\[3\] u_cpu.rf_ram.memory\[93\]\[3\] u_cpu.rf_ram.memory\[94\]\[3\]
+ u_cpu.rf_ram.memory\[95\]\[3\] _02075_ _01847_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09240__I _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__A1 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06361_ _01515_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11606__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08100_ u_cpu.rf_ram.memory\[74\]\[5\] _03416_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09080_ u_cpu.rf_ram.memory\[131\]\[7\] _04038_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08651__A1 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06292_ u_cpu.rf_ram.memory\[96\]\[2\] u_cpu.rf_ram.memory\[97\]\[2\] u_cpu.rf_ram.memory\[98\]\[2\]
+ u_cpu.rf_ram.memory\[99\]\[2\] _01938_ _01824_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08031_ u_cpu.rf_ram.memory\[129\]\[4\] _03376_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11538__A1 u_cpu.rf_ram.memory\[89\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11756__CLK net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A1 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09982_ _04629_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__A2 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06104__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08933_ _02984_ _03550_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08706__A2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08864_ _03647_ _03903_ _03912_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06568__I1 u_cpu.rf_ram.memory\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05943__I _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07815_ u_cpu.rf_ram.memory\[48\]\[7\] _03211_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06812__S1 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08795_ u_cpu.rf_ram.memory\[71\]\[4\] _03868_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07746_ _03182_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10277__B2 _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ _02914_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07142__A1 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09416_ _04251_ _04267_ _04270_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06628_ _01724_ _02271_ _01702_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08890__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10029__A1 _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09150__I _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10029__B2 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09347_ _04165_ _04217_ _04223_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06559_ u_cpu.rf_ram.memory\[20\]\[5\] u_cpu.rf_ram.memory\[21\]\[5\] u_cpu.rf_ram.memory\[22\]\[5\]
+ u_cpu.rf_ram.memory\[23\]\[5\] _01891_ _02003_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12531__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06328__S0 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10229__C _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09278_ _04180_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08229_ _03343_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06723__B _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11240_ _05570_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09198__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12681__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10201__A1 _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08945__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11171_ _05525_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10752__A2 _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10122_ _04801_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06014__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10053_ _04694_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10504__A2 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06559__I1 u_cpu.rf_ram.memory\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05853__I _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06803__S1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__A1 _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ _05317_ _05388_ _05393_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11629__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07133__A1 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10886_ _05350_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08881__A1 u_cpu.rf_ram.memory\[138\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06731__I1 u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12625_ _01122_ net266 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__S0 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08633__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _01054_ net313 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11779__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11507_ u_cpu.rf_ram.memory\[100\]\[1\] _05743_ _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12487_ _00988_ net242 u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09189__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11438_ u_cpu.rf_ram.memory\[25\]\[6\] _05698_ _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06247__I0 u_cpu.rf_ram.memory\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ _01449_ _04236_ _04233_ _02499_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10743__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout396_I net397 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06262__I3 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _01546_ _01557_ _01566_ _01575_ _01578_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13039_ u_scanchain_local.data_out net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12404__CLK net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__A2 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05861_ u_cpu.cpu.csr_imm u_cpu.rf_ram_if.rtrig0 _01456_ _01464_ _01510_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_39_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _03034_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05792_ u_cpu.cpu.decode.opcode\[2\] _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__A1 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07531_ _03038_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12554__CLK net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07462_ _02971_ _02987_ _02992_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07675__A2 _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ _04127_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06413_ _02055_ _02057_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07393_ _02881_ u_cpu.rf_ram_if.wdata0_r\[5\] _02936_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_143_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ _03537_ _03454_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06344_ _01758_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08624__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07427__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06486__I0 u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ _04038_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06275_ u_cpu.rf_ram.memory\[56\]\[2\] u_cpu.rf_ram.memory\[57\]\[2\] u_cpu.rf_ram.memory\[58\]\[2\]
+ u_cpu.rf_ram.memory\[59\]\[2\] _01623_ _01812_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08014_ _03350_ _03359_ _03367_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10065__B _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09965_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _04604_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08916_ u_cpu.rf_ram.memory\[137\]\[0\] _03947_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09896_ u_cpu.rf_ram.memory\[113\]\[4\] _04589_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12084__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10498__A1 _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09352__A2 _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _03901_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07363__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06166__A2 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06797__S0 _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07902__A3 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ u_cpu.rf_ram.memory\[73\]\[6\] _03851_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ u_cpu.rf_ram.memory\[51\]\[1\] _03171_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07115__A1 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10740_ u_cpu.rf_ram.memory\[97\]\[1\] _05260_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08863__A1 u_cpu.rf_ram.memory\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11921__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _05204_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12410_ _00911_ net485 u_cpu.rf_ram.memory\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07418__A2 _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11997__D _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12341_ _00842_ net350 u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08091__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10973__A2 _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05848__I _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12272_ _00773_ net255 u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11223_ _05562_ _05552_ _05563_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ u_cpu.rf_ram.memory\[84\]\[3\] _05518_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09591__A2 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _04772_ _04775_ _04786_ _04787_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11085_ _05469_ _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10036_ _04667_ _04696_ _04723_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06788__S0 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12577__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08894__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07106__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11987_ _00509_ net223 u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06628__B _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08854__A1 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10938_ u_cpu.rf_ram.memory\[103\]\[4\] _05380_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07657__A2 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__B1 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10110__C2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10661__A1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout144_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10869_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _05341_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06180__I2 u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12608_ _01105_ net447 u_cpu.rf_ram.memory\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout311_I net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12539_ _01040_ net328 u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout409_I net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10964__A2 _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06093__A1 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06060_ _01705_ _01708_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05840__A1 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09031__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__A2 _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout408 net409 net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout419 net421 net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_98_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07593__A1 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06396__A2 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09750_ _04236_ _02611_ u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.mem_bytecnt\[0\] _04482_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06962_ _02474_ u_cpu.rf_ram.rdata\[5\] _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05913_ _01551_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08701_ _03806_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09681_ _04170_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06893_ _02524_ _02521_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11141__A2 _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _03647_ _03759_ _03768_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05844_ _01476_ _01485_ _01490_ _01494_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06699__A3 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11944__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08563_ _03666_ _03718_ _03721_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ _03025_ _03015_ _03026_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07648__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _03352_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout15 net16 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout26 net27 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10652__A1 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07445_ _02944_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout37 net38 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout48 net51 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout59 net60 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06320__A2 _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07376_ u_cpu.rf_ram.memory\[82\]\[2\] _02922_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ _04070_ _04065_ _04072_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10404__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06327_ _01971_ _01973_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08073__A2 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09270__A1 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07281__B1 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09046_ _03993_ _04027_ _04029_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06258_ _01560_ _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05831__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09022__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06189_ _01607_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07883__I _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09573__A2 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11380__A2 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _03274_ u_arbiter.i_wb_cpu_rdt\[8\] _04639_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09879_ _02690_ _04574_ _04581_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11132__A2 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11910_ _00432_ net275 u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12890_ _01387_ net507 u_cpu.rf_ram.memory\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07887__A2 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10891__A1 _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11841_ _00363_ net98 u_cpu.rf_ram.memory\[67\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08219__I _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11772_ _00294_ net91 u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__I _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10643__A1 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10723_ _02871_ _05233_ _04949_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10654_ _04077_ _05185_ _05192_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11199__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08064__A2 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10585_ _05149_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06183__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12324_ _00825_ net468 u_cpu.rf_ram.memory\[34\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05822__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12255_ _00756_ net349 u_cpu.rf_ram.memory\[38\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11817__CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10159__B1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11206_ _05512_ _02961_ _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09564__A2 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12186_ _00700_ net373 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ u_cpu.rf_ram.memory\[69\]\[5\] _05505_ _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11967__CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05976__I2 u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11068_ _05411_ _05457_ _05464_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11123__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10019_ _03274_ u_arbiter.i_wb_cpu_rdt\[14\] _04707_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_3_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10659__I _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout261_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout359_I net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10634__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout526_I net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06302__A2 _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ _02609_ u_scanchain_local.module_data_in\[56\] _02796_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06805__C _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07161_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _02727_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_34_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08055__A2 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10937__A2 _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__C _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06112_ u_cpu.rf_ram.memory\[128\]\[0\] u_cpu.rf_ram.memory\[129\]\[0\] u_cpu.rf_ram.memory\[130\]\[0\]
+ u_cpu.rf_ram.memory\[131\]\[0\] _01759_ _01760_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07092_ _02629_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06456__I3 u_cpu.rf_ram.memory\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05813__A1 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06043_ _01498_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout205 net206 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06369__A2 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout216 net228 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11362__A2 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout227 net228 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09802_ u_arbiter.i_wb_cpu_rdt\[6\] _04512_ _04524_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xfanout238 net239 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07994_ _03353_ _03331_ _03354_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout249 net251 net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10570__B1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09733_ u_cpu.rf_ram.memory\[33\]\[0\] _04472_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06945_ _02582_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11114__A2 _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07869__A2 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09664_ _04427_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06876_ _02513_ _02515_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05951__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08615_ _03757_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05827_ u_cpu.cpu.immdec.imm24_20\[1\] _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09595_ _04346_ _04378_ _04385_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06541__A2 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08546_ _03668_ _03706_ _03711_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08818__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10625__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _03666_ _03663_ _03667_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09491__A1 _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ _02954_ _02966_ _02968_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12272__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ _02907_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11050__A1 u_cpu.rf_ram.memory\[106\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _04228_ _02874_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06152__S1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09029_ _04014_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12040_ _00554_ net25 u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06604__I0 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12942_ u_cpu.cpu.o_wdata0 net336 u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10700__C _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12873_ _01370_ net501 u_cpu.rf_ram.memory\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06178__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11824_ _00346_ net203 u_cpu.rf_ram.memory\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12615__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10616__A1 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__A2 _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11755_ _00277_ net393 u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__I2 u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06296__A1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10706_ _05223_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11686_ _00208_ net464 u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06391__S1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10637_ u_cpu.rf_ram.memory\[3\]\[7\] _05171_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09234__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12765__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07096__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07245__B1 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10568_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _05137_ _05139_ _02800_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06143__S1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12307_ _00808_ net196 u_cpu.rf_ram.memory\[92\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10499_ u_cpu.rf_ram.memory\[30\]\[1\] _05096_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout107_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08412__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12238_ _00013_ net281 u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07548__A1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12169_ _00683_ net80 u_cpu.rf_ram.memory\[130\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout476_I net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12145__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06730_ _01476_ _02323_ _02372_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput5 io_in[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09243__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06661_ u_cpu.rf_ram.memory\[36\]\[6\] u_cpu.rf_ram.memory\[37\]\[6\] u_cpu.rf_ram.memory\[38\]\[6\]
+ u_cpu.rf_ram.memory\[39\]\[6\] _01679_ _01680_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_92_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08400_ u_cpu.rf_ram.memory\[19\]\[2\] _03613_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09380_ _04234_ u_cpu.cpu.state.o_cnt_r\[2\] _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12295__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06592_ _01692_ _02207_ _02216_ _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_80_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10607__A1 u_cpu.rf_ram.memory\[109\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _03568_ _03565_ _03569_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10458__I1 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A2 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08262_ _03525_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10083__A2 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06382__S1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07213_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _02779_ _02781_ _02703_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08028__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09225__A1 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _03440_ _03480_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07144_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07087__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06107__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07075_ _02674_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06551__B _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05946__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06026_ u_cpu.rf_ram.memory\[120\]\[0\] u_cpu.rf_ram.memory\[121\]\[0\] u_cpu.rf_ram.memory\[122\]\[0\]
+ u_cpu.rf_ram.memory\[123\]\[0\] _01673_ _01674_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06211__B2 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ u_cpu.rf_ram.memory\[40\]\[3\] _03338_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11099__A1 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09716_ _04431_ _04459_ _04462_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06928_ _02557_ _02518_ _02558_ _02566_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_60_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09153__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12638__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09700__A2 _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09647_ _04337_ _04414_ _04417_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06859_ u_cpu.cpu.decode.op22 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07711__A1 u_cpu.rf_ram.memory\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ u_cpu.rf_ram.memory\[118\]\[7\] _04364_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ u_cpu.rf_ram.memory\[55\]\[4\] _03698_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09464__A1 u_cpu.rf_ram.memory\[92\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11662__CLK net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08267__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12788__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06278__A1 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11540_ u_cpu.rf_ram.memory\[89\]\[7\] _05753_ _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07401__I _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__S1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _02971_ _05718_ _05723_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08019__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__A1 _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11023__A1 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10422_ _05051_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07078__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12018__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07778__A1 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10231__C1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10762__I _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ u_cpu.cpu.immdec.imm19_12_20\[7\] _04947_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05856__I u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07049__S _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09519__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08232__I _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06450__B2 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _04942_ _04943_ _04944_ _04601_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12168__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12023_ _00537_ net43 u_cpu.rf_ram.memory\[140\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10711__B _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07950__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09063__I _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12925_ _01422_ net384 u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06505__A2 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12856_ _01353_ net334 u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11807_ _00329_ net127 u_cpu.rf_ram.memory\[76\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09455__A1 u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08258__A2 _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12787_ _01284_ net108 u_cpu.rf_ram.memory\[84\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11262__A1 _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11738_ _00260_ net288 u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout224_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10873__S _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11669_ _00191_ net463 u_cpu.rf_ram.memory\[45\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11014__A1 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11565__A2 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10672__I _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__A2 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07900_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _03287_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ _03857_ _03915_ _03922_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07831_ u_cpu.rf_ram.memory\[47\]\[4\] _03237_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09930__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07941__A1 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__I2 u_cpu.rf_ram.memory\[98\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ _03146_ _03186_ _03193_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09501_ _04253_ _04321_ _04326_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10828__A1 u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06713_ u_cpu.rf_ram.memory\[72\]\[6\] u_cpu.rf_ram.memory\[73\]\[6\] u_cpu.rf_ram.memory\[74\]\[6\]
+ u_cpu.rf_ram.memory\[75\]\[6\] _01694_ _01695_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07693_ _02945_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11685__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09694__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08497__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12930__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06644_ _01523_ _02286_ _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06052__S0 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09432_ _03271_ _04229_ _04278_ _04279_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06575_ u_cpu.rf_ram.memory\[32\]\[5\] u_cpu.rf_ram.memory\[33\]\[5\] u_cpu.rf_ram.memory\[34\]\[5\]
+ u_cpu.rf_ram.memory\[35\]\[5\] _01745_ _02024_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09363_ u_cpu.cpu.mem_bytecnt\[0\] _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08249__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11253__A1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08314_ _03503_ _03552_ _03558_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09294_ u_cpu.rf_ram.memory\[123\]\[7\] _04180_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _03493_ _03514_ _03516_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06680__A1 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11005__A1 _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09749__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _03408_ _03469_ _03471_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11556__A2 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07127_ _02709_ _02710_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12310__CLK net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07058_ _02664_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11308__A2 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06009_ _01656_ _01657_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06983__A2 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12460__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07932__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06586__I2 u_cpu.rf_ram.memory\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10819__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06300__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _05399_ _05401_ _05403_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12710_ _01207_ net151 u_cpu.rf_ram.memory\[104\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11492__A1 u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10757__I _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12641_ _01138_ net143 u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11362__B _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09437__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11244__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__A2 _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12572_ _01070_ net323 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07131__I _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11523_ _05753_ _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__A2 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06510__I2 u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06671__A1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11454_ u_cpu.rf_ram.memory\[24\]\[4\] _05710_ _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11547__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10405_ u_cpu.rf_ram.memory\[31\]\[4\] _05039_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11385_ u_cpu.rf_ram.memory\[27\]\[0\] _05671_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06191__B _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10336_ _04963_ _04965_ _04636_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12803__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06974__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ u_cpu.cpu.immdec.imm7 _02851_ _04884_ _04928_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08176__A1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12006_ _00520_ net45 u_cpu.rf_ram.memory\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10198_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _04773_ _04866_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07923__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06210__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout174_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09676__A1 u_cpu.rf_ram.memory\[122\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12908_ _01405_ net200 u_cpu.rf_ram.memory\[98\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10286__A2 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09521__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10667__I _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout341_I net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12839_ _01336_ net118 u_cpu.rf_ram.memory\[87\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout439_I net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06360_ _01512_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10038__A2 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09979__A2 _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06291_ _01548_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07976__I _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ _03341_ _03372_ _03378_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06662__A1 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11538__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09600__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _04660_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ _03943_ _03947_ _03956_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout87_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ u_cpu.rf_ram.memory\[14\]\[7\] _03901_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07814_ _02951_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06273__S0 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08794_ _03853_ _03864_ _03870_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07390__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07745_ _02957_ _03100_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09667__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07676_ _03129_ _03134_ _03136_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ u_cpu.rf_ram.memory\[90\]\[1\] _04268_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09419__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06627_ u_cpu.rf_ram.memory\[76\]\[5\] u_cpu.rf_ram.memory\[77\]\[5\] u_cpu.rf_ram.memory\[78\]\[5\]
+ u_cpu.rf_ram.memory\[79\]\[5\] _01979_ _01726_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06740__I2 u_cpu.rf_ram.memory\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11226__A1 _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10029__A2 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06558_ _01719_ _02201_ _02001_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09346_ u_cpu.rf_ram.memory\[36\]\[3\] _04221_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06328__S1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06489_ _01599_ _02133_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09277_ _04180_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08642__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07886__I _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06653__A1 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _03503_ _03495_ _03504_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12826__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ _03456_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10201__A2 _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11170_ _05473_ _05526_ _05529_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _04801_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06956__A2 u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12976__CLK net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08158__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__I1 u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _02493_ _04699_ _04738_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06708__A2 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06559__I2 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06264__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12206__CLK net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06030__I _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09658__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ u_cpu.rf_ram.memory\[104\]\[2\] _05392_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12356__CLK net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ _02960_ _05158_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08881__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11217__A1 _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06892__A1 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12624_ _01121_ net263 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12555_ _00023_ net313 u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08633__A2 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11506_ _03620_ _05742_ _05744_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12486_ _00987_ net242 u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _05632_ _05695_ _05702_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08397__A1 u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11368_ u_cpu.cpu.genblk3.csr.mie_mtie _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10319_ _04733_ _04727_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_45_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11299_ _05555_ _05607_ _05610_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08149__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08420__I _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13038_ net536 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout291_I net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout389_I net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09897__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13038__I net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05860_ _01500_ _01508_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__A1 u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ u_cpu.cpu.decode.co_mem_word u_cpu.cpu.bne_or_bge u_cpu.cpu.csr_d_sel _01442_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_94_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _03038_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06875__I _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08321__A1 u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07461_ u_cpu.rf_ram.memory\[81\]\[2\] _02991_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06412_ _01483_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09200_ _04127_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07392_ _02876_ u_cpu.rf_ram_if.wdata1_r\[5\] _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11723__CLK net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06343_ u_cpu.rf_ram.memory\[128\]\[2\] u_cpu.rf_ram.memory\[129\]\[2\] u_cpu.rf_ram.memory\[130\]\[2\]
+ u_cpu.rf_ram.memory\[131\]\[2\] _01759_ _01760_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09131_ _03729_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06824__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06635__A1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ _03166_ _04013_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06274_ _01919_ _01920_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10346__B _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08013_ u_cpu.rf_ram.memory\[119\]\[6\] _03362_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11873__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11021__I _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06115__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06399__B1 _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06938__A2 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _04604_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08915_ _03945_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09895_ _04436_ _04585_ _04591_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09888__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08846_ _03901_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10498__A2 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06797__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08777_ _03751_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05989_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ _03129_ _03170_ _03172_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08312__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07115__A2 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ _03023_ _03118_ _03124_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06174__I0 u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10670_ _02918_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09329_ _04168_ _04205_ _04212_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06734__B _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06626__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12340_ _00841_ net479 u_cpu.rf_ram.memory\[120\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13004__CLK net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12271_ _00772_ net359 u_cpu.rf_ram.memory\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11222_ u_cpu.rf_ram.memory\[85\]\[4\] _05558_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06025__I _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10186__A1 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A2 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11153_ _05475_ _05514_ _05519_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05864__I _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _04680_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11084_ _05204_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_1_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09879__A1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10035_ _02617_ _04720_ _04722_ _04683_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_48_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08551__A1 u_cpu.rf_ram.memory\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06788__S1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11986_ _00508_ net214 u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _05320_ _05376_ _05382_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10110__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__A2 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__B2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10010__I _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10661__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10868_ _05330_ _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_34_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12607_ _01104_ net447 u_cpu.rf_ram.memory\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06180__I3 u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_83_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11896__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10799_ _05196_ _05295_ _05297_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06617__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10413__A2 _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12538_ _01039_ net328 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10166__B _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10881__S _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__A1 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout304_I net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12469_ _00970_ net491 u_cpu.rf_ram.memory\[114\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05840__A2 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09031__A2 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10680__I _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout409 net451 net409 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09246__I _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07593__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08150__I _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06961_ _02584_ _02593_ _02594_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ _03736_ _03807_ _03810_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05912_ _01503_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_100_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12521__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06228__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09680_ _04438_ _04428_ _04439_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06892_ u_cpu.cpu.bufreg.lsb\[0\] _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08542__A1 u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08631_ u_cpu.rf_ram.memory\[9\]\[7\] _03757_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05843_ _01493_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ u_cpu.rf_ram.memory\[53\]\[1\] _03719_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09098__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12671__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07513_ u_cpu.rf_ram.memory\[20\]\[4\] _03021_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10101__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08493_ _03677_ _03664_ _03678_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11016__I _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout16 net20 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06856__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout27 net32 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10652__A2 _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07444_ _02978_ _02967_ _02979_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout38 net40 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net51 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07375_ _02900_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13027__CLK net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06554__B _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05949__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09114_ u_cpu.rf_ram.memory\[12\]\[2\] _04071_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10404__A2 _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06326_ u_cpu.rf_ram.memory\[64\]\[2\] u_cpu.rf_ram.memory\[65\]\[2\] u_cpu.rf_ram.memory\[66\]\[2\]
+ u_cpu.rf_ram.memory\[67\]\[2\] _01720_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08325__I _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06257_ u_cpu.rf_ram.memory\[8\]\[2\] u_cpu.rf_ram.memory\[9\]\[2\] u_cpu.rf_ram.memory\[10\]\[2\]
+ u_cpu.rf_ram.memory\[11\]\[2\] _01561_ _01564_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07281__A1 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09045_ u_cpu.rf_ram.memory\[132\]\[0\] _04028_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05831__A2 _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ _01659_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__A2 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11619__CLK net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__I _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08781__A1 u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09947_ _02705_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08995__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ u_arbiter.i_wb_cpu_rdt\[29\] _04511_ _04497_ u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08533__A1 u_cpu.rf_ram.memory\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08829_ u_cpu.rf_ram.memory\[143\]\[1\] _03890_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10340__A1 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11840_ _00362_ net98 u_cpu.rf_ram.memory\[67\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10891__A2 _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11771_ _00293_ net91 u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ _02870_ _02618_ _02873_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10643__A2 _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06162__I3 u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10653_ u_cpu.rf_ram.memory\[2\]\[5\] _05188_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08235__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _02832_ _05144_ _05146_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09261__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12323_ _00824_ net487 u_cpu.rf_ram.memory\[34\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05822__A2 _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12254_ _00755_ net349 u_cpu.rf_ram.memory\[38\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10159__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09013__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10159__B2 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10714__B _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11205_ _05195_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12544__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__S0 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12185_ _00699_ net372 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _05480_ _05501_ _05508_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11067_ u_cpu.rf_ram.memory\[107\]\[4\] _05461_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10018_ _04604_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06639__B _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout254_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11969_ _00491_ net31 u_cpu.rf_ram.memory\[53\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10634__A2 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout421_I net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10675__I _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout519_I net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__12074__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06111_ _01721_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07263__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__I _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06042_ _01494_ _01666_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout206 net229 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout217 net219 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _04526_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08763__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout228 net229 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07993_ u_cpu.rf_ram.memory\[40\]\[7\] _03329_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout239 net244 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _04470_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06944_ _02484_ _02556_ _02567_ _02581_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_45_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09663_ _03101_ _04426_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10322__A1 _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06875_ _02514_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08614_ _03757_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05826_ u_cpu.cpu.immdec.imm19_12_20\[5\] u_cpu.rf_ram_if.rtrig0 _01477_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06621__S0 _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09594_ u_cpu.rf_ram.memory\[121\]\[5\] _04381_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07224__I u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06541__A3 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ u_cpu.rf_ram.memory\[54\]\[2\] _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08818__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10625__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12417__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ u_cpu.rf_ram.memory\[57\]\[1\] _03664_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09491__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ u_cpu.rf_ram.memory\[21\]\[0\] _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07358_ _02906_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10389__A1 u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ _01949_ _01951_ _01953_ _01955_ _01689_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_104_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06301__I0 u_cpu.rf_ram.memory\[124\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _02843_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09028_ _03998_ _04015_ _04018_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08754__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__A1 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12941_ u_cpu.rf_ram_if.wdata0_r\[6\] net336 u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10313__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06612__S0 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12872_ _01369_ net500 u_cpu.rf_ram.memory\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11823_ _00345_ net203 u_cpu.rf_ram.memory\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08809__A2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__B1 _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06973__I _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12097__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11754_ _00276_ net429 u_cpu.rf_ram.memory\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09482__A2 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07070__S _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _04677_ _05231_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11685_ _00207_ net374 u_cpu.rf_ram.memory\[51\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10636_ _04079_ _05173_ _05181_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09234__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__A2 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07245__A1 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07245__B2 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _05109_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12306_ _00807_ net198 u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07796__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11934__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10498_ _04800_ _05095_ _05097_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12237_ _00012_ net279 u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10163__C _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12168_ _00682_ net84 u_cpu.rf_ram.memory\[130\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11119_ u_cpu.rf_ram.memory\[108\]\[6\] _05493_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12099_ _00613_ net264 u_cpu.rf_ram.memory\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout371_I net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout469_I net470 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09170__A1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06660_ _02296_ _02298_ _02300_ _02302_ _01740_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07181__B1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06591_ _01795_ _02225_ _02234_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_91_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07979__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ u_cpu.rf_ram.memory\[62\]\[1\] _03566_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06816__C _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07484__A1 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ _03068_ _03087_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02752_ _02780_
+ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08192_ _03166_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09225__A2 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06039__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11032__A2 _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07143_ _02704_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07087__I1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__A3 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08984__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07074_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_dbus_dat\[18\] _02671_ _02674_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10791__A1 u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ _01607_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07539__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06123__I _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07976_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05962__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09434__I _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09715_ u_cpu.rf_ram.memory\[116\]\[1\] _04460_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06927_ _02562_ _02565_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09646_ u_cpu.rf_ram.memory\[112\]\[1\] _04415_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06858_ u_cpu.cpu.state.o_cnt_r\[3\] _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05809_ _01443_ _01444_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09577_ _04348_ _04366_ _04374_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06789_ _01615_ _02430_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11807__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08528_ _03671_ _03694_ _03700_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__I3 u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06278__A2 _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11271__A2 _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08459_ u_cpu.rf_ram.memory\[58\]\[3\] _03654_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11470_ u_cpu.rf_ram.memory\[0\]\[2\] _05722_ _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11957__CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09216__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07227__A1 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10421_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _05048_
+ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11023__A2 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10231__B1 _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10231__C2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10352_ u_cpu.cpu.immdec.imm19_12_20\[8\] _04698_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10283_ u_cpu.cpu.immdec.imm7 _02462_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12022_ _00536_ net43 u_cpu.rf_ram.memory\[140\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__I _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05872__I _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07065__S _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09152__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12924_ _01421_ net383 u_cpu.rf_ram.memory\[89\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12855_ _01352_ net286 u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12732__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07799__I _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11806_ _00328_ net128 u_cpu.rf_ram.memory\[76\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12786_ _01283_ net112 u_cpu.rf_ram.memory\[84\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07466__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11262__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11737_ _00259_ net288 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11668_ _00190_ net461 u_cpu.rf_ram.memory\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09207__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12882__CLK net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10619_ _03037_ _03480_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10953__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout217_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11599_ _00121_ net414 u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07769__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08966__A1 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10773__A1 u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__A2 _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06292__I2 u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07830_ _03220_ _03233_ _03239_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06878__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12262__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ u_cpu.rf_ram.memory\[41\]\[5\] _03189_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09500_ u_cpu.rf_ram.memory\[34\]\[2\] _04325_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09143__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06712_ _01711_ _02354_ _01715_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07692_ _03146_ _03135_ _03147_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07154__B1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09694__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06347__I3 u_cpu.rf_ram.memory\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09431_ _03273_ _04242_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06643_ u_cpu.rf_ram.memory\[28\]\[6\] u_cpu.rf_ram.memory\[29\]\[6\] u_cpu.rf_ram.memory\[30\]\[6\]
+ u_cpu.rf_ram.memory\[31\]\[6\] _01524_ _01525_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06052__S1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06901__B1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09362_ _03271_ _04231_ _04232_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_fanout32_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06574_ _01796_ _02217_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__I _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ u_cpu.rf_ram.memory\[63\]\[3\] _03556_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07457__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06504__I0 u_cpu.rf_ram.memory\[100\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11253__A2 _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09293_ _04174_ _04182_ _04190_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08244_ u_cpu.rf_ram.memory\[65\]\[0\] _03515_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11005__A2 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ u_cpu.rf_ram.memory\[68\]\[0\] _03470_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__B _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05957__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08957__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07126_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08333__I _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10764__A1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07057_ _02608_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08709__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06008_ u_cpu.rf_ram.memory\[108\]\[0\] u_cpu.rf_ram.memory\[109\]\[0\] u_cpu.rf_ram.memory\[110\]\[0\]
+ u_cpu.rf_ram.memory\[111\]\[0\] _01549_ _01563_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12605__CLK net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__A2 _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07932__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06586__I3 u_cpu.rf_ram.memory\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ _03011_ _03100_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_25_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ u_cpu.rf_ram.memory\[99\]\[0\] _05402_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09685__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ u_cpu.rf_ram.memory\[11\]\[2\] _04406_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11492__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12640_ _01137_ net143 u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11244__A2 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12571_ _01069_ net327 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11522_ _02898_ _03182_ _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06510__I3 u_cpu.rf_ram.memory\[107\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12135__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11453_ _05628_ _05706_ _05712_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05867__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__A1 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _04810_ _05035_ _05041_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08243__I _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11384_ _05669_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10755__A1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__A1 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10335_ _04765_ _04823_ _04964_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12285__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10266_ _04925_ _04926_ _04927_ _02851_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10507__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09373__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12005_ _00519_ net45 u_cpu.rf_ram.memory\[142\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08176__A2 _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06187__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10197_ _04616_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09676__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12907_ _01404_ net200 u_cpu.rf_ram.memory\[98\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10948__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout167_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12838_ _01335_ net111 u_cpu.rf_ram.memory\[87\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10169__B _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12769_ _01266_ net138 u_cpu.rf_ram.memory\[108\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout334_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06290_ _01511_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10994__A1 _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout501_I net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10683__I _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06662__A2 _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__A1 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08153__I _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12628__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10746__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09600__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07611__A1 u_cpu.rf_ram.memory\[78\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _04601_ _04669_ _04671_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ u_cpu.rf_ram.memory\[137\]\[7\] _03945_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12778__CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ _03644_ _03903_ _03911_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06178__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ _03226_ _03213_ _03227_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08793_ u_cpu.rf_ram.memory\[71\]\[3\] _03868_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06273__S1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07744_ _03103_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07678__A1 u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11474__A2 _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07675_ u_cpu.rf_ram.memory\[45\]\[0\] _03135_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09414_ _04246_ _04267_ _04269_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06626_ _01705_ _02269_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09419__A2 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06740__I3 u_cpu.rf_ram.memory\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ _04161_ _04217_ _04222_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06557_ u_cpu.rf_ram.memory\[24\]\[5\] u_cpu.rf_ram.memory\[25\]\[5\] u_cpu.rf_ram.memory\[26\]\[5\]
+ u_cpu.rf_ram.memory\[27\]\[5\] _01746_ _01774_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11226__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06102__A1 _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09276_ _03196_ _04179_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06488_ u_cpu.rf_ram.memory\[40\]\[4\] u_cpu.rf_ram.memory\[41\]\[4\] u_cpu.rf_ram.memory\[42\]\[4\]
+ u_cpu.rf_ram.memory\[43\]\[4\] _02027_ _01601_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08227_ u_cpu.rf_ram.memory\[66\]\[3\] _03501_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06653__A2 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07850__A1 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _02915_ _03457_ _03460_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ _02628_ _02623_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06405__A2 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08089_ _03336_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10120_ _02890_ _04426_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__A2 _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09355__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06008__I2 u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10051_ _04720_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06311__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06264__S1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A1 u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11465__A2 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _05387_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__A2 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10884_ _05349_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12623_ _01120_ net263 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__11217__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06892__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12554_ _00024_ net313 u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11505_ u_cpu.rf_ram.memory\[100\]\[0\] _05743_ _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06644__A2 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12485_ _00986_ net243 u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06495__I2 u_cpu.rf_ram.memory\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09069__I _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09969__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11436_ u_cpu.rf_ram.memory\[25\]\[5\] _05698_ _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11367_ _05657_ _05638_ _05658_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10318_ _04645_ _04687_ _04790_ _04821_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__I _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11298_ u_cpu.rf_ram.memory\[87\]\[1\] _05608_ _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09346__A1 u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _04909_ _04911_ _04824_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11153__A1 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09897__A2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10879__S _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout284_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10900__A1 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05790_ u_cpu.cpu.immdec.imm24_20\[0\] _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06580__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09649__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout451_I net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11456__A2 _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07460_ _02986_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ u_cpu.rf_ram.memory\[104\]\[3\] u_cpu.rf_ram.memory\[105\]\[3\] u_cpu.rf_ram.memory\[106\]\[3\]
+ u_cpu.rf_ram.memory\[107\]\[3\] _02056_ _01571_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06722__I3 u_cpu.rf_ram.memory\[135\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07391_ _02901_ _02934_ _02935_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__I _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09130_ _04081_ _04066_ _04082_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06342_ _01752_ _01988_ _01756_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08085__A1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10967__A1 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06824__C _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _04011_ _04028_ _04037_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07832__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06635__A2 _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06273_ u_cpu.rf_ram.memory\[60\]\[2\] u_cpu.rf_ram.memory\[61\]\[2\] u_cpu.rf_ram.memory\[62\]\[2\]
+ u_cpu.rf_ram.memory\[63\]\[2\] _01617_ _01619_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08012_ _03347_ _03359_ _03366_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10719__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08388__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06399__B2 _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09963_ _04613_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08914_ _03945_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09894_ u_cpu.rf_ram.memory\[113\]\[3\] _04589_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11144__A1 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09888__A2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08845_ _03900_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07899__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08560__A2 _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ _03857_ _03846_ _03858_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06571__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05970__I _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05988_ _01591_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07727_ u_cpu.rf_ram.memory\[51\]\[0\] _03171_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11447__A2 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ u_cpu.rf_ram.memory\[46\]\[3\] _03122_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06323__B2 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06609_ _01604_ _02252_ _01640_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07589_ _03025_ _03070_ _03077_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ u_cpu.rf_ram.memory\[37\]\[4\] _04209_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__A1 u_cpu.rf_ram.memory\[77\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07823__A1 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _02931_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12455__D _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06182__S0 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12943__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12270_ _00771_ net359 u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11221_ _05211_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10186__A2 _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11152_ u_cpu.rf_ram.memory\[84\]\[2\] _05518_ _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10103_ _04776_ _04778_ _04785_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11083_ _05473_ _05470_ _05474_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09879__A2 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10034_ _04721_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__A1 u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12323__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05880__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11438__A2 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11985_ _00507_ net214 u_cpu.rf_ram.memory\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05813__C _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A2 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10936_ u_cpu.rf_ram.memory\[103\]\[3\] _05380_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12473__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__I3 u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10867_ _05340_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12606_ _01103_ net443 u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ u_cpu.rf_ram.memory\[96\]\[0\] _05296_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10949__A1 u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06617__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12537_ _01038_ net328 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12468_ _00969_ net491 u_cpu.rf_ram.memory\[114\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06093__A3 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11419_ _05634_ _05683_ _05691_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12399_ _00900_ net454 u_cpu.rf_ram.memory\[116\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10182__B _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout499_I net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09319__A1 u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06960_ _02583_ u_cpu.rf_ram_if.rdata1\[4\] _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ _01559_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06228__S1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06891_ _02520_ _02526_ _02529_ u_cpu.cpu.state.stage_two_req _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_45_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _03644_ _03759_ _03767_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08542__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05842_ _01491_ _01492_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__I u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12816__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ _03661_ _03718_ _03720_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07512_ _02933_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ u_cpu.rf_ram.memory\[57\]\[6\] _03669_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10101__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout17 net20 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07443_ u_cpu.rf_ram.memory\[21\]\[5\] _02972_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout28 net30 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout39 net40 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11840__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12966__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08058__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ _02920_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08606__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ _04064_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout9_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06325_ _01517_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09044_ _04026_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06256_ _01785_ _01901_ _01902_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06126__I _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__A1 u_cpu.rf_ram.memory\[120\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06187_ _01667_ _01834_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10168__A2 _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12346__CLK net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08781__A2 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _04634_ _04635_ _04636_ _04637_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_132_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _04579_ _04580_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09730__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08828_ _03843_ _03889_ _03891_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12496__CLK net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ u_cpu.rf_ram.memory\[73\]\[0\] _03846_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11207__I _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08297__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11770_ _00292_ net393 u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10721_ _05238_ _05244_ _05246_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08049__A1 u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ _04075_ _05184_ _05191_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10267__B _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07420__I _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10583_ _05148_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06155__S0 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12322_ _00823_ net467 u_cpu.rf_ram.memory\[34\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06036__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09549__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12253_ _00754_ net348 u_cpu.rf_ram.memory\[38\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10159__A2 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05875__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11204_ _02982_ _05540_ _05549_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08221__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12184_ _00698_ net372 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06458__S1 _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08772__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ u_cpu.rf_ram.memory\[69\]\[4\] _05505_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11713__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12839__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11066_ _05409_ _05457_ _05463_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10730__B _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09721__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _02706_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11863__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12989__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11968_ _00490_ net30 u_cpu.rf_ram.memory\[53\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09810__I _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A1 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ u_cpu.rf_ram.memory\[102\]\[5\] _05367_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06838__A2 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout247_I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11899_ _00421_ net372 u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12219__CLK net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09788__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout414_I net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06110_ _01541_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07090_ _02682_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08460__A1 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12369__CLK net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10691__I _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06041_ _01671_ _01677_ _01682_ _01688_ _01689_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__11347__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08212__A1 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout207 net208 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09800_ _04497_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09960__A1 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout218 net219 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout229 net230 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07992_ _03352_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10570__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09731_ _04470_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06943_ _02518_ _02532_ _02554_ _02580_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09662_ _03355_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06874_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01462_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06526__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07505__I _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10322__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08613_ _03037_ _03183_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_94_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09921__S _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05825_ _01470_ _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09593_ _04344_ _04377_ _04384_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06621__S1 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08544_ _03705_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06129__I1 u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06829__A2 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08475_ _03333_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07426_ _02965_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10881__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__I _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10087__B _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _02905_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06308_ _01683_ _01954_ _01687_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07288_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _02843_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ u_cpu.rf_ram.memory\[133\]\[1\] _04016_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06239_ u_cpu.rf_ram.memory\[28\]\[2\] u_cpu.rf_ram.memory\[29\]\[2\] u_cpu.rf_ram.memory\[30\]\[2\]
+ u_cpu.rf_ram.memory\[31\]\[2\] _01504_ _01771_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11736__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__A1 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06765__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09929_ _04605_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09703__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11886__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12940_ u_cpu.rf_ram_if.wdata0_r\[5\] net336 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11510__A1 u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10313__A2 _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12871_ _01368_ net498 u_cpu.rf_ram.memory\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06612__S1 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11822_ _00344_ net203 u_cpu.rf_ram.memory\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10077__A1 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10776__I _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11753_ _00275_ net429 u_cpu.rf_ram.memory\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__B2 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _05226_ _05229_ _05230_ _04776_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11684_ _00206_ net374 u_cpu.rf_ram.memory\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10635_ u_cpu.rf_ram.memory\[3\]\[6\] _05176_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10566_ _05138_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10725__B _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12305_ _00806_ net198 u_cpu.rf_ram.memory\[92\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10497_ u_cpu.rf_ram.memory\[30\]\[0\] _05096_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12236_ _00011_ net280 u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12661__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09942__A1 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08745__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12167_ _00681_ net79 u_cpu.rf_ram.memory\[130\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06756__A1 _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11118_ _05482_ _05490_ _05497_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12098_ _00612_ net344 u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout197_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13017__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11049_ _05413_ _05445_ _05452_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11501__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__A2 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12041__CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06590_ _02227_ _02229_ _02231_ _02233_ _01489_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout531_I net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11609__CLK net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _03511_ _03515_ _03524_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07211_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\] u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__12191__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08191_ _03426_ _03470_ _03479_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ _02714_ _02720_ _02723_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10240__A1 _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07073_ _02673_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06995__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10791__A2 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ _01605_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06047__I0 u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ _02926_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09714_ _04425_ _04459_ _04461_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06926_ _01442_ _02563_ _02564_ _02548_ _02549_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_95_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09645_ _04332_ _04414_ _04416_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06857_ _01447_ _01450_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _01447_ _01450_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09576_ u_cpu.rf_ram.memory\[118\]\[6\] _04369_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06788_ u_cpu.rf_ram.memory\[92\]\[7\] u_cpu.rf_ram.memory\[93\]\[7\] u_cpu.rf_ram.memory\[94\]\[7\]
+ u_cpu.rf_ram.memory\[95\]\[7\] _02075_ _01619_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10059__A1 _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ u_cpu.rf_ram.memory\[55\]\[3\] _03698_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__S0 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12534__CLK net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08458_ _03570_ _03650_ _03655_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07409_ _02950_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ _03579_ _03598_ _03606_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11559__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10420_ _05050_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _04600_ _05001_ _05003_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_87_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06986__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06314__I _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10282_ _02869_ _02534_ _04674_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12021_ _00535_ net45 u_cpu.rf_ram.memory\[140\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08727__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10534__A2 _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07145__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09152__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12923_ _01420_ net383 u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10298__B2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06597__S0 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06984__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12854_ _01351_ net286 u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06910__A1 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07081__S _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _00327_ net127 u_cpu.rf_ram.memory\[76\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12785_ _01282_ net112 u_cpu.rf_ram.memory\[84\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08663__A1 _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11736_ _00258_ net337 u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11667_ _00189_ net461 u_cpu.rf_ram.memory\[45\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10618_ _04818_ _05161_ _05170_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11598_ _00120_ net414 u_cpu.rf_ram.memory\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10222__A1 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06277__I0 u_cpu.rf_ram.memory\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout112_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10549_ _05128_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06977__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11130__I _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10773__A2 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12219_ _00733_ net348 u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12407__CLK net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout481_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07760_ _03144_ _03185_ _03192_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09143__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06711_ u_cpu.rf_ram.memory\[68\]\[6\] u_cpu.rf_ram.memory\[69\]\[6\] u_cpu.rf_ram.memory\[70\]\[6\]
+ u_cpu.rf_ram.memory\[71\]\[6\] _01712_ _01713_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07691_ u_cpu.rf_ram.memory\[45\]\[5\] _03140_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07154__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06588__S0 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _02614_ _02616_ _02613_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_65_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06642_ _01476_ _02236_ _02285_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06901__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06901__B2 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _02498_ u_cpu.cpu.state.o_cnt\[2\] _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_94_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06573_ u_cpu.rf_ram.memory\[36\]\[5\] u_cpu.rf_ram.memory\[37\]\[5\] u_cpu.rf_ram.memory\[38\]\[5\]
+ u_cpu.rf_ram.memory\[39\]\[5\] _01797_ _01680_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08312_ _03500_ _03552_ _03557_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08654__A1 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09292_ u_cpu.rf_ram.memory\[123\]\[6\] _04185_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout25_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06504__I1 u_cpu.rf_ram.memory\[101\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08243_ _03513_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06760__S0 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08614__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08174_ _03468_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08406__A1 u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06680__A3 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10213__A1 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07125_ _02708_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10764__A2 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06134__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07056_ _02663_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06007_ _01628_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09906__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08709__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05973__I _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06196__A2 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07393__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07958_ _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06909_ u_cpu.cpu.state.o_cnt_r\[0\] _02501_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07889_ _03277_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09628_ _04401_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08893__A1 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11924__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ _04350_ _04354_ _04363_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11215__I _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12570_ _01068_ net323 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08645__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11521_ _03646_ _05743_ _05752_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06751__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11452_ u_cpu.rf_ram.memory\[24\]\[3\] _05710_ _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08524__I _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__I0 u_cpu.rf_ram.memory\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10403_ u_cpu.rf_ram.memory\[31\]\[3\] _05039_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10204__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11383_ _05669_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10755__A2 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06044__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _04596_ _02642_ _04987_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10265_ _02534_ _04926_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10507__A2 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__S _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12004_ _00518_ net56 u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09373__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ _04862_ _04673_ _04863_ _04722_ _04780_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06026__I3 u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07384__A1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06187__A2 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11180__A2 _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout390 net391 net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07136__A1 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12906_ _01403_ net205 u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08884__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12837_ _01334_ net101 u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11125__I _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06219__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12768_ _01265_ net138 u_cpu.rf_ram.memory\[108\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11719_ _00241_ net387 u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout327_I net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12699_ _01196_ net136 u_cpu.rf_ram.memory\[102\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06742__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10994__A2 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08434__I _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09061__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10746__A2 _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ _03941_ _03947_ _03955_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ u_cpu.rf_ram.memory\[14\]\[6\] _03906_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06178__A2 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07812_ u_cpu.rf_ram.memory\[48\]\[6\] _03218_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08792_ _03850_ _03864_ _03869_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11947__CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _03150_ _03171_ _03180_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07127__A1 _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ _03133_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07678__A2 _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08875__A1 u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08609__I _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10682__A1 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09413_ u_cpu.rf_ram.memory\[90\]\[0\] _04268_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06625_ u_cpu.rf_ram.memory\[72\]\[5\] u_cpu.rf_ram.memory\[73\]\[5\] u_cpu.rf_ram.memory\[74\]\[5\]
+ u_cpu.rf_ram.memory\[75\]\[5\] _01867_ _01695_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11035__I _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06350__A2 _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08627__A1 u_cpu.rf_ram.memory\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06556_ _01523_ _02199_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09344_ u_cpu.rf_ram.memory\[36\]\[2\] _04221_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09275_ _03355_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06487_ _01559_ _02131_ _01801_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06102__A2 _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06733__S0 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05968__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ _03340_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07850__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08157_ u_cpu.rf_ram.memory\[6\]\[1\] _03458_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05861__B2 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07108_ _02630_ u_scanchain_local.module_data_in\[37\] _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _03413_ _03410_ _03414_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07039_ _02654_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06661__I0 u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _04724_ _04725_ _04727_ _04728_ _04736_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__I3 u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11162__A2 _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12872__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10952_ _05315_ _05388_ _05391_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08519__I _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__I _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10883_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _05330_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12622_ _01119_ net263 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08618__A1 u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12553_ _01053_ net184 u_cpu.rf_ram.memory\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08094__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09291__A1 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06724__S0 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11504_ _05741_ _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12484_ _00985_ net242 u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11435_ _05630_ _05694_ _05701_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11366_ u_cpu.cpu.genblk3.csr.mstatus_mie _05638_ _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09594__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06247__I3 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _04865_ _04971_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11297_ _05550_ _05607_ _05609_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09346__A2 _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10248_ _04826_ _04910_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10024__I _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _04847_ _04843_ _04848_ _04799_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout277_I net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08857__A1 u_cpu.rf_ram.memory\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08429__I _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout444_I net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ _01605_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07390_ u_cpu.rf_ram.memory\[82\]\[4\] _02922_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06341_ u_cpu.rf_ram.memory\[140\]\[2\] u_cpu.rf_ram.memory\[141\]\[2\] u_cpu.rf_ram.memory\[142\]\[2\]
+ u_cpu.rf_ram.memory\[143\]\[2\] _01753_ _01754_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08085__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10967__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09060_ u_cpu.rf_ram.memory\[132\]\[7\] _04026_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06272_ _01581_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06486__I3 u_cpu.rf_ram.memory\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08011_ u_cpu.rf_ram.memory\[119\]\[5\] _03362_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07596__A1 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06399__A2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11392__A2 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06643__I0 u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _04650_ _04653_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06412__I _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08913_ _03182_ _03887_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12895__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09893_ _04433_ _04585_ _04590_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07348__A1 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11144__A2 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08844_ _03256_ _03083_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07899__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05987_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08775_ u_cpu.rf_ram.memory\[73\]\[5\] _03851_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07726_ _03169_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08848__A1 u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08339__I _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07657_ _03020_ _03118_ _03123_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09879__B _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06323__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07520__A1 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06174__I2 u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06608_ u_cpu.rf_ram.memory\[116\]\[5\] u_cpu.rf_ram.memory\[117\]\[5\] u_cpu.rf_ram.memory\[118\]\[5\]
+ u_cpu.rf_ram.memory\[119\]\[5\] _02069_ _01638_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07588_ u_cpu.rf_ram.memory\[80\]\[4\] _03074_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12275__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06539_ _01724_ _02183_ _01738_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09327_ _04165_ _04205_ _04211_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08076__A2 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09273__A1 u_cpu.rf_ram.memory\[124\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06706__S0 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__A1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07284__B1 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _04165_ _04154_ _04166_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07823__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06182__S1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08209_ u_cpu.rf_ram.memory\[67\]\[6\] _03486_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10109__I _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09189_ u_cpu.rf_ram.memory\[127\]\[3\] _04120_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11220_ _05560_ _05552_ _05561_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07587__A1 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _05513_ _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10102_ _04684_ _04780_ _04784_ _04660_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09328__A2 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11082_ u_cpu.rf_ram.memory\[83\]\[1\] _05471_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10033_ _04656_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08000__A2 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10894__A1 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A2 _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11984_ _00506_ net221 u_cpu.rf_ram.memory\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12618__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06197__C _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09500__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10935_ _05317_ _05376_ _05381_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07511__A1 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06165__I2 u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10866_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _05335_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10728__B _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12605_ _01102_ net443 u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12768__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11642__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11403__I _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10797_ _05294_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11071__A1 u_cpu.rf_ram.memory\[107\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12536_ _01037_ net330 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05825__A1 _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12467_ _00968_ net491 u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06941__B _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ u_cpu.rf_ram.memory\[26\]\[6\] _05686_ _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11792__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12398_ _00899_ net458 u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06660__C _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11374__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06625__I0 u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10421__I1 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11349_ _05641_ _05645_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10582__B1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12148__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout394_I net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11126__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ _01558_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13019_ _00080_ net533 u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06890_ _01452_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _02528_ u_cpu.cpu.state.init_done
+ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_66_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10885__A1 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05841_ u_cpu.cpu.immdec.imm24_20\[3\] _01473_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07750__A1 u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06553__A2 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08159__I _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08560_ u_cpu.rf_ram.memory\[53\]\[0\] _03719_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_2_540 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_66_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07511_ _03023_ _03015_ _03024_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08491_ _03349_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07442_ _02938_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout18 net20 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout29 net30 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ _02919_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08058__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11313__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09112_ _02920_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06324_ _01704_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06069__B2 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09043_ _04026_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06255_ _01533_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__A2 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ u_cpu.rf_ram.memory\[124\]\[1\] u_cpu.rf_ram.memory\[125\]\[1\] u_cpu.rf_ram.memory\[126\]\[1\]
+ u_cpu.rf_ram.memory\[127\]\[1\] _01668_ _01669_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07569__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08230__A2 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09945_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _04603_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11117__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09876_ u_arbiter.i_wb_cpu_rdt\[28\] _04495_ _04519_ u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05981__I _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09730__A2 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ u_cpu.rf_ram.memory\[143\]\[0\] _03890_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06298__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06395__I2 u_cpu.rf_ram.memory\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _03844_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10628__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ u_cpu.rf_ram.memory\[44\]\[2\] _03159_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A2 _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _03749_ _03796_ _03803_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12910__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10720_ _02871_ _05233_ _05245_ _04787_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ u_cpu.rf_ram.memory\[2\]\[4\] _05188_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08049__A2 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11053__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _05144_ _05146_ _02832_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06155__S1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05807__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12321_ _00822_ net487 u_cpu.rf_ram.memory\[34\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__B _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09549__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12252_ _00753_ net339 u_cpu.rf_ram.memory\[38\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11356__A2 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11203_ u_cpu.rf_ram.memory\[10\]\[7\] _05538_ _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12183_ _00697_ net373 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08221__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11134_ _05478_ _05501_ _05507_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11108__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A2 _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11065_ u_cpu.rf_ram.memory\[107\]\[3\] _05461_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05891__I _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10730__C _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09363__I u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10016_ _04640_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07732__A1 u_cpu.rf_ram.memory\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06535__A2 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10619__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09485__A1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11967_ _00489_ net30 u_cpu.rf_ram.memory\[53\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12590__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11292__A1 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A2 _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10918_ _05322_ _05363_ _05370_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11898_ _00420_ net372 u_cpu.rf_ram.memory\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout142_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10849_ _03276_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_32_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11044__A1 u_cpu.rf_ram.memory\[106\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06227__I _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10972__I _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12519_ _01020_ net311 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout407_I net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06471__A1 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06040_ _01488_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__I _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08212__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07058__I _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net211 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout219 net227 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07991_ _02950_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09730_ _02984_ _03130_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06942_ _00798_ _02572_ _02579_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ _04151_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06873_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11688__CLK net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10322__A3 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08612_ _03755_ _03733_ _03756_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12933__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05824_ _01472_ _01474_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_54_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ u_cpu.rf_ram.memory\[121\]\[4\] _04381_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08543_ _03666_ _03706_ _03709_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09476__A1 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08279__A2 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06129__I2 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08474_ _03661_ _03663_ _03665_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07521__I _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06385__S1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07425_ _02965_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06137__I _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07356_ u_cpu.rf_ram_if.wdata0_r\[0\] _02902_ _02904_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_52_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06307_ u_cpu.rf_ram.memory\[116\]\[2\] u_cpu.rf_ram.memory\[117\]\[2\] u_cpu.rf_ram.memory\[118\]\[2\]
+ u_cpu.rf_ram.memory\[119\]\[2\] _01684_ _01685_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07287_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _02826_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06238_ _01497_ _01821_ _01885_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _03993_ _04015_ _04017_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05896__S0 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08352__I _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ u_cpu.rf_ram.memory\[48\]\[1\] u_cpu.rf_ram.memory\[49\]\[1\] u_cpu.rf_ram.memory\[50\]\[1\]
+ u_cpu.rf_ram.memory\[51\]\[1\] _01636_ _01638_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09400__A1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08203__A2 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10546__B1 _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12463__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__A2 _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _04619_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09703__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09859_ u_arbiter.i_wb_cpu_rdt\[22\] _04559_ _04560_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__I2 u_cpu.rf_ram.memory\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07714__A1 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11218__I _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11510__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10122__I _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06073__S0 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12870_ _01367_ net496 u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09911__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11821_ _00343_ net203 u_cpu.rf_ram.memory\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__A1 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06756__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__A2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11752_ _00274_ net429 u_cpu.rf_ram.memory\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__S1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _04672_ _04714_ _04865_ _04891_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09219__A1 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11683_ _00205_ net391 u_cpu.rf_ram.memory\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08690__A2 _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10634_ _04077_ _05173_ _05180_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09786__C _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10565_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _05137_ _05132_ u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _00805_ net198 u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08262__I _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10496_ _05094_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12235_ _00010_ net287 u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12166_ _00680_ net80 u_cpu.rf_ram.memory\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07953__A1 u_cpu.rf_ram.memory\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11117_ u_cpu.rf_ram.memory\[108\]\[5\] _05493_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12956__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12097_ _00611_ net343 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11048_ u_cpu.rf_ram.memory\[106\]\[5\] _05448_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07705__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10032__I _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11980__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09458__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout357_I net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12999_ _00058_ net526 u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08437__I _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout524_I net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07210_ _02778_ _02775_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08190_ u_cpu.rf_ram.memory\[68\]\[7\] _03468_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07141_ _02721_ u_scanchain_local.module_data_in\[41\] _02722_ u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09630__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06295__I1 u_cpu.rf_ram.memory\[109\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10240__A2 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_dbus_dat\[17\] _02671_ _02673_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12486__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06023_ _01659_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06995__A2 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08197__A1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07974_ _03337_ _03330_ _03339_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09713_ u_cpu.rf_ram.memory\[116\]\[0\] _04460_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06420__I _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06925_ _02485_ _02522_ u_cpu.cpu.alu.cmp_r _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09644_ u_cpu.rf_ram.memory\[112\]\[0\] _04415_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06856_ _02495_ _02489_ _02493_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10700__B1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05807_ u_cpu.cpu.decode.op21 _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _04346_ _04366_ _04373_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06787_ _01580_ _02419_ _02428_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_71_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10059__A2 _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08526_ _03668_ _03694_ _03699_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08121__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__S1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ u_cpu.rf_ram.memory\[58\]\[2\] _03654_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08672__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ _02949_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08388_ u_cpu.rf_ram.memory\[60\]\[6\] _03601_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12829__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11559__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07339_ _02887_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08082__I _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _02715_ _02646_ _04739_ _05002_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06986__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09009_ _03745_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10281_ _04835_ _04759_ _04940_ _04941_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12979__CLK net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12020_ _00534_ net61 u_cpu.rf_ram.memory\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08810__I _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__A1 u_cpu.rf_ram.memory\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06738__A2 _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11495__A1 _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12922_ _01419_ net383 u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__A1 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12853_ _01350_ net286 u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12359__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06910__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11247__A1 u_cpu.rf_ram.memory\[110\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11804_ _00326_ net127 u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12784_ _01281_ net112 u_cpu.rf_ram.memory\[84\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11735_ _00257_ net285 u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08663__A2 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11666_ _00188_ net462 u_cpu.rf_ram.memory\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10617_ u_cpu.rf_ram.memory\[109\]\[7\] _05159_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09612__A1 u_cpu.rf_ram.memory\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11597_ _00119_ net189 u_cpu.rf_ram.memory\[81\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10222__A2 _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _02758_ _05123_ _05125_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06977__A2 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout105_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10479_ _05082_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12218_ _00732_ net300 u_cpu.rf_ram.memory\[125\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09915__A2 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07926__A1 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06729__A2 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _00663_ net52 u_cpu.rf_ram.memory\[132\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout474_I net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06710_ _01971_ _02352_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06037__S0 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11486__A1 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ _02939_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__A1 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__S1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06641_ _02275_ _02284_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11238__A1 u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ _02498_ u_cpu.cpu.state.o_cnt\[2\] _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06572_ _02209_ _02211_ _02213_ _02215_ _01740_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_94_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08311_ u_cpu.rf_ram.memory\[63\]\[2\] _03556_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _04171_ _04182_ _04189_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08654__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08242_ _03513_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout18_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11876__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08173_ _03468_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09603__A1 u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08406__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10213__A2 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07124_ _02707_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07055_ u_arbiter.i_wb_cpu_rdt\[13\] u_arbiter.i_wb_cpu_dbus_dat\[10\] _02658_ _02663_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06006_ _01651_ _01653_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09906__A2 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07917__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07957_ _02906_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11477__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06908_ _02531_ _02533_ _02538_ _02546_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ _03275_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _03276_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06579__S1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ _04068_ _04402_ _04405_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ u_cpu.cpu.alu.i_rs1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11229__A1 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09558_ u_cpu.rf_ram.memory\[120\]\[7\] _04352_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12651__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ u_cpu.rf_ram.memory\[56\]\[4\] _03686_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _04262_ _04310_ _04318_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06200__S0 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11520_ u_cpu.rf_ram.memory\[100\]\[7\] _05741_ _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__I _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__S1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11451_ _05625_ _05706_ _05711_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06408__A1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10402_ _04807_ _05035_ _05040_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11401__A1 _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__I _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__A2 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11382_ _05310_ _03196_ _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09070__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _04596_ u_arbiter.i_wb_cpu_rdt\[17\] _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _02614_ _04281_ u_cpu.cpu.decode.opcode\[1\] _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07908__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12003_ _00517_ net56 u_cpu.rf_ram.memory\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10195_ _04712_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07384__A2 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout380 net381 net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__12181__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout391 net392 net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11468__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12905_ _01402_ net203 u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10140__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06195__I0 u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08884__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12836_ _01333_ net101 u_cpu.rf_ram.memory\[87\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12767_ _01264_ net136 u_cpu.rf_ram.memory\[108\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11899__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11718_ _00240_ net387 u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08715__I _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12698_ _01195_ net136 u_cpu.rf_ram.memory\[102\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06742__S1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout222_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11649_ _00171_ net395 u_cpu.rf_ram.memory\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09061__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12524__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08860_ _03641_ _03903_ _03910_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08572__A1 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07811_ _02945_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ u_cpu.rf_ram.memory\[71\]\[2\] _03868_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11459__A1 _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07742_ u_cpu.rf_ram.memory\[51\]\[7\] _03169_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10421__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__A1 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07673_ _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10131__A1 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06186__I0 u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08875__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11316__I _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09412_ _04266_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06430__S0 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06886__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06624_ _01862_ _02267_ _01865_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10682__A2 _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09343_ _04216_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06555_ u_cpu.rf_ram.memory\[28\]\[5\] u_cpu.rf_ram.memory\[29\]\[5\] u_cpu.rf_ram.memory\[30\]\[5\]
+ u_cpu.rf_ram.memory\[31\]\[5\] _01524_ _01771_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08627__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09274_ _04177_ _04155_ _04178_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06486_ u_cpu.rf_ram.memory\[32\]\[4\] u_cpu.rf_ram.memory\[33\]\[4\] u_cpu.rf_ram.memory\[34\]\[4\]
+ u_cpu.rf_ram.memory\[35\]\[4\] _01745_ _02024_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06733__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08225_ _03500_ _03495_ _03502_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ _02908_ _03457_ _03459_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05861__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09052__A2 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ _02692_ _02643_ _02693_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06497__S0 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ u_cpu.rf_ram.memory\[74\]\[1\] _03411_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07038_ u_arbiter.i_wb_cpu_rdt\[5\] u_arbiter.i_wb_cpu_dbus_dat\[2\] _02652_ _02654_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08563__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__A1 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ u_cpu.rf_ram.memory\[135\]\[6\] _03986_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08315__A1 u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06748__C _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ u_cpu.rf_ram.memory\[104\]\[1\] _05389_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06877__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10673__A2 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05924__I0 u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10882_ _05348_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12621_ _01118_ net263 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08618__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12552_ _01052_ net188 u_cpu.rf_ram.memory\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10286__B _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06483__C _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11503_ _05741_ _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06724__S1 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12483_ _00984_ net241 u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11434_ u_cpu.rf_ram.memory\[25\]\[4\] _05698_ _05701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06055__I _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10189__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06488__S0 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11365_ u_cpu.cpu.genblk3.csr.mstatus_mpie _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05894__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07087__S _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10316_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _04773_ _04971_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11296_ u_cpu.rf_ram.memory\[87\]\[0\] _05608_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10247_ _04724_ _04753_ _04822_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08554__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10361__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10178_ u_cpu.cpu.immdec.imm24_20\[3\] _04841_ _04674_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07109__A2 _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout172_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10113__A1 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08857__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06868__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__A2 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__I _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12819_ _01316_ net125 u_cpu.rf_ram.memory\[110\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout437_I net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06340_ _01469_ _01986_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08445__I _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09282__A2 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06715__S1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06271_ _01910_ _01912_ _01914_ _01917_ _01613_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_15_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09985__B _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08010_ _03344_ _03358_ _03365_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06479__S0 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07596__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11914__CLK net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _04652_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _03943_ _03928_ _03944_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09892_ u_cpu.rf_ram.memory\[113\]\[2\] _04589_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03861_ _03890_ _03899_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ _03748_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05986_ _01501_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07524__I u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07725_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08848__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10655__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ u_cpu.rf_ram.memory\[46\]\[2\] _03122_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__A2 _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06607_ _02065_ _02250_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ _03023_ _03070_ _03076_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05979__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__A2 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ u_cpu.rf_ram.memory\[37\]\[3\] _04209_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ u_cpu.rf_ram.memory\[76\]\[4\] u_cpu.rf_ram.memory\[77\]\[4\] u_cpu.rf_ram.memory\[78\]\[4\]
+ u_cpu.rf_ram.memory\[79\]\[4\] _01979_ _01726_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_16_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09273__A2 _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06706__S1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07284__A1 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__A2 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ u_cpu.rf_ram.memory\[124\]\[3\] _04162_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06469_ _01513_ _02113_ _02001_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08208_ _03422_ _03483_ _03490_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09025__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _04090_ _04116_ _04121_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08139_ u_cpu.rf_ram.memory\[75\]\[3\] _03446_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11594__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A2 _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11150_ _05473_ _05514_ _05517_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08090__I _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10101_ _04650_ _04781_ _04783_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10125__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11081_ _05201_ _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08536__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _04680_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10343__A1 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10061__S _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10894__A2 _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11983_ _00505_ net421 u_cpu.rf_ram.memory\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10934_ u_cpu.rf_ram.memory\[103\]\[2\] _05380_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07511__A2 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10865_ _05339_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06570__I0 u_cpu.rf_ram.memory\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05889__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12604_ _01101_ net442 u_cpu.rf_ram.memory\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _05294_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12535_ _01036_ net330 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05825__A2 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12466_ _00967_ net490 u_cpu.rf_ram.memory\[114\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11937__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09016__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06941__C _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11417_ _05632_ _05683_ _05690_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12397_ _00898_ net458 u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11348_ _03273_ _05642_ _05644_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11279_ _05555_ _05595_ _05598_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13018_ _00079_ net533 u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10334__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout387_I net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05840_ u_cpu.cpu.immdec.imm19_12_20\[7\] _01471_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10885__A2 _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_2_541 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07510_ u_cpu.rf_ram.memory\[20\]\[3\] _03021_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _03675_ _03664_ _03676_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ _02976_ _02966_ _02977_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06561__I0 u_cpu.rf_ram.memory\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout19 net20 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_62_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12712__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _02918_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ _04068_ _04065_ _04069_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06323_ _01960_ _01964_ _01967_ _01969_ _01858_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _03012_ _04013_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06254_ u_cpu.rf_ram.memory\[0\]\[2\] u_cpu.rf_ram.memory\[1\]\[2\] u_cpu.rf_ram.memory\[2\]\[2\]
+ u_cpu.rf_ram.memory\[3\]\[2\] _01786_ _01900_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12862__CLK net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07018__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06185_ _01823_ _01826_ _01829_ _01831_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06616__I1 u_cpu.rf_ram.memory\[81\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06423__I _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06777__B1 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _02726_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ u_arbiter.i_wb_cpu_dbus_dat\[28\] _04521_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10325__A1 _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _03888_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12242__CLK net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08757_ _03844_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05969_ _01551_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ _03154_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10628__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ u_cpu.rf_ram.memory\[141\]\[5\] _03799_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07639_ _03023_ _03106_ _03112_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05930__C _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12392__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11504__I _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10650_ _04073_ _05184_ _05190_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ _04168_ _04193_ _04200_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11053__A2 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10581_ _05147_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _00821_ net488 u_cpu.rf_ram.memory\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09909__I _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10261__B1 _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10800__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07009__A1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12251_ _00752_ net339 u_cpu.rf_ram.memory\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11202_ _02980_ _05540_ _05548_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07429__I _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12182_ _00696_ net372 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11133_ u_cpu.rf_ram.memory\[69\]\[3\] _05505_ _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _05406_ _05457_ _05462_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10015_ _04703_ _04635_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12735__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10619__A2 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11966_ _00488_ net30 u_cpu.rf_ram.memory\[53\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09485__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10917_ u_cpu.rf_ram.memory\[102\]\[4\] _05367_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11897_ _00419_ net270 u_cpu.rf_ram.memory\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10848_ _05328_ _05313_ _05329_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout135_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10779_ _05196_ _05283_ _05285_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12518_ _01019_ net311 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12115__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12449_ _00950_ net482 u_cpu.rf_ram.memory\[113\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout302_I net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08748__A1 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06243__I _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout209 net211 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07990_ _03350_ _03331_ _03351_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12265__CLK net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06941_ _02577_ _02578_ _01463_ _02510_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10307__A1 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__A1 u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06606__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _04350_ _04415_ _04424_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06872_ _02484_ _02511_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08611_ u_cpu.rf_ram.memory\[52\]\[7\] _03731_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05823_ u_cpu.cpu.immdec.imm24_20\[4\] _01473_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09591_ _04342_ _04377_ _04383_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06782__I0 u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08542_ u_cpu.rf_ram.memory\[54\]\[1\] _03707_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout48_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__I _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09476__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08473_ u_cpu.rf_ram.memory\[57\]\[0\] _03664_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ _02961_ _02964_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__A2 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07355_ u_cpu.rf_ram_if.wdata1_r\[0\] _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06306_ _01678_ _01952_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08987__A1 u_cpu.rf_ram.memory\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__C2 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06837__I1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ _02701_ u_scanchain_local.module_data_in\[67\] _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10794__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06581__C _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09025_ u_cpu.rf_ram.memory\[133\]\[0\] _04016_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06237_ _01874_ _01884_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06462__A2 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05896__S1 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__A1 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12608__CLK net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06153__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06168_ _01629_ _01815_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09400__A2 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10546__B2 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07411__A1 u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06099_ _01637_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _04612_ _04618_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11632__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12758__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09858_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _04557_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07714__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08911__A1 u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06073__S1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08809_ _03848_ _03876_ _03879_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09789_ _04490_ _04516_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _00342_ net199 u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11751_ _00273_ net430 u_cpu.rf_ram.memory\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06525__I0 u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11234__I _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _04776_ _05228_ _04739_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10278__C _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11682_ _00204_ net389 u_cpu.rf_ram.memory\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09219__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10633_ u_cpu.rf_ram.memory\[3\]\[5\] _05176_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11026__A2 _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12138__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06772__B _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10234__B1 _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08978__A1 u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10564_ _05106_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10294__B _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06989__B1 _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12303_ _00804_ net198 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10495_ _05094_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12288__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06063__I _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12234_ _00009_ net285 u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12165_ _00679_ net79 u_cpu.rf_ram.memory\[130\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07953__A2 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11116_ _05480_ _05489_ _05496_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12096_ _00610_ net338 u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11409__I _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09155__A1 _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11047_ _05411_ _05444_ _05451_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07705__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08902__A1 u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12998_ _00057_ net525 u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11265__A2 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout252_I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11949_ _00471_ net27 u_cpu.rf_ram.memory\[55\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10188__C _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11017__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout517_I net518 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10076__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08969__A1 u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07140_ _02624_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07641__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07071_ _02672_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06295__I2 u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07069__I _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06022_ _01667_ _01670_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11655__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09394__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08197__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12900__CLK net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07973_ u_cpu.rf_ram.memory\[40\]\[2\] _03338_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11319__I _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09146__A1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09712_ _04458_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06924_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02479_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_64_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09643_ _04413_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06855_ _02485_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__I0 u_cpu.rf_ram.memory\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10700__A1 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10700__B2 _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05806_ u_cpu.cpu.decode.op26 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ u_cpu.rf_ram.memory\[118\]\[5\] _04369_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06380__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06786_ _02421_ _02423_ _02425_ _02427_ _02072_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_97_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__A2 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08525_ u_cpu.rf_ram.memory\[55\]\[2\] _03698_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11256__A2 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11054__I _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08121__A2 _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06148__I _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08456_ _03649_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07407_ _02948_ _02582_ _02881_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07880__A1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _03577_ _03598_ _03605_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05987__I _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07338_ u_cpu.raddr\[0\] _02886_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12430__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A2 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07269_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _02828_ _02713_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _04003_ _03995_ _04004_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10280_ _04599_ _04681_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08188__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12580__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07935__A2 _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09688__A2 _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12921_ _01418_ net382 u_cpu.rf_ram.memory\[89\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06746__I0 u_cpu.rf_ram.memory\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__A2 _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12852_ _01349_ net334 u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08538__I _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07442__I _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _00325_ net165 u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12783_ _01280_ net118 u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12000__D _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08112__A2 _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06058__I _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11734_ _00256_ net316 u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11665_ _00187_ net461 u_cpu.rf_ram.memory\[45\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10616_ _04816_ _05161_ _05169_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _00118_ net215 u_cpu.rf_ram.memory\[81\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11678__CLK net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ _05127_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07623__A1 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ u_arbiter.i_wb_cpu_dbus_adr\[30\] u_arbiter.i_wb_cpu_dbus_adr\[31\] _05078_
+ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09376__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12217_ _00731_ net343 u_cpu.rf_ram.memory\[125\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11183__A1 _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12148_ _00662_ net53 u_cpu.rf_ram.memory\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10930__A1 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12079_ _00593_ net227 u_cpu.rf_ram.memory\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06037__S1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout467_I net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06737__I0 u_cpu.rf_ram.memory\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12303__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08351__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06640_ _02277_ _02279_ _02281_ _02283_ _01470_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_25_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06571_ _01468_ _02214_ _01792_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09300__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08103__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03551_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09290_ u_cpu.rf_ram.memory\[123\]\[5\] _04185_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10997__A1 u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _02985_ _03087_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10419__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07301__B _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ _03013_ _03087_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09603__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07123_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__A1 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11410__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07054_ _02662_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06005_ _01595_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07917__A2 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09943__S _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10921__A1 u_cpu.rf_ram.memory\[102\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07956_ _03228_ _03315_ _03324_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06907_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02545_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11477__A2 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07887_ u_arbiter.i_wb_cpu_ack _02702_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09626_ u_cpu.rf_ram.memory\[11\]\[1\] _04403_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06838_ _02465_ _02478_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08358__I _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11229__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09557_ _04348_ _04354_ _04362_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06769_ u_cpu.rf_ram.memory\[100\]\[7\] u_cpu.rf_ram.memory\[101\]\[7\] u_cpu.rf_ram.memory\[102\]\[7\]
+ u_cpu.rf_ram.memory\[103\]\[7\] _01569_ _01543_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _03671_ _03682_ _03688_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ u_cpu.rf_ram.memory\[35\]\[6\] _04313_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08439_ u_cpu.rf_ram.memory\[5\]\[5\] _03632_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06200__S1 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12946__CLK net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11450_ u_cpu.rf_ram.memory\[24\]\[2\] _05710_ _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08093__I _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ u_cpu.rf_ram.memory\[31\]\[2\] _05039_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06259__I2 u_cpu.rf_ram.memory\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11401__A2 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10128__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__A3 _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11381_ _03271_ u_cpu.cpu.genblk3.csr.timer_irq_r _05021_ _05668_ _01358_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ u_cpu.cpu.immdec.imm19_12_20\[6\] _04970_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11970__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09358__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10263_ u_cpu.cpu.immdec.imm19_12_20\[0\] _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12002_ _00007_ net283 u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08030__A1 _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10194_ _04703_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06592__A1 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout370 net371 net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout381 net384 net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout392 net397 net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11468__A2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09530__A1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12904_ _01401_ net205 u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08268__I _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06195__I1 u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10140__A2 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12835_ _01332_ net129 u_cpu.rf_ram.memory\[111\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12766_ _01263_ net138 u_cpu.rf_ram.memory\[108\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11717_ _00239_ net402 u_cpu.rf_ram.memory\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12697_ _01194_ net136 u_cpu.rf_ram.memory\[102\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11648_ _00170_ net395 u_cpu.rf_ram.memory\[42\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09597__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11579_ _00101_ net210 u_cpu.rf_ram.memory\[82\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout215_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09827__I _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09349__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _03224_ _03213_ _03225_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08572__A2 _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ _03863_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06583__A1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07741_ _03148_ _03171_ _03179_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12819__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11459__A2 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ _03130_ _03132_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10131__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ _04266_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06623_ u_cpu.rf_ram.memory\[68\]\[5\] u_cpu.rf_ram.memory\[69\]\[5\] u_cpu.rf_ram.memory\[70\]\[5\]
+ u_cpu.rf_ram.memory\[71\]\[5\] _01712_ _01863_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06430__S1 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06886__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _04158_ _04217_ _04220_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06554_ _01497_ _02148_ _02198_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout30_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09273_ u_cpu.rf_ram.memory\[124\]\[7\] _04153_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06485_ _01796_ _02129_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11332__I _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ u_cpu.rf_ram.memory\[66\]\[2\] _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06426__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11993__CLK net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ u_cpu.rf_ram.memory\[6\]\[0\] _03458_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11395__A1 _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07106_ _02684_ u_scanchain_local.module_data_in\[36\] _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08086_ _03333_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08260__A1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06497__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12349__CLK net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ _02653_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12499__CLK net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08988_ _03939_ _03983_ _03990_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10370__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07939_ _03313_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08315__A2 _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ _05309_ _05388_ _05390_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _04070_ _04389_ _04394_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06421__S1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10881_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _05330_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12620_ _01117_ net148 u_cpu.rf_ram.memory\[93\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08079__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12551_ _01051_ net188 u_cpu.rf_ram.memory\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11502_ _03012_ _05157_ _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12482_ _00983_ net239 u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09579__A1 _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11433_ _05628_ _05694_ _05700_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11386__A1 _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10189__A2 _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11364_ _05656_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06488__S1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10315_ _04952_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06652__I2 u_cpu.rf_ram.memory\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11295_ _05606_ _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11138__A1 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11716__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10246_ _04908_ _04673_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08003__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09751__A1 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08554__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__I2 u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ u_cpu.cpu.immdec.imm24_20\[2\] _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06565__A1 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09382__I _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09503__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08306__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06317__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11310__A1 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06868__A2 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout165_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12818_ _01315_ net131 u_cpu.rf_ram.memory\[110\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout332_I net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12749_ _01246_ net115 u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10196__C _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06270_ _01915_ _01916_ _01807_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08490__A1 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10991__I _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06479__S1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08793__A2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _02707_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _04651_ _04652_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11129__A1 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08911_ u_cpu.rf_ram.memory\[39\]\[7\] _03926_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09891_ _04584_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10432__S _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ u_cpu.rf_ram.memory\[143\]\[7\] _03888_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10352__A2 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07805__I _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _03855_ _03845_ _03856_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05985_ _01598_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07724_ _03166_ _03168_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12791__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07655_ _03117_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06606_ u_cpu.rf_ram.memory\[112\]\[5\] u_cpu.rf_ram.memory\[113\]\[5\] u_cpu.rf_ram.memory\[114\]\[5\]
+ u_cpu.rf_ram.memory\[115\]\[5\] _02066_ _01840_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07586_ u_cpu.rf_ram.memory\[80\]\[3\] _03074_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12021__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _04161_ _04205_ _04210_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06537_ _01705_ _02181_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11062__I _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06167__S0 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09256_ _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06468_ u_cpu.rf_ram.memory\[24\]\[4\] u_cpu.rf_ram.memory\[25\]\[4\] u_cpu.rf_ram.memory\[26\]\[4\]
+ u_cpu.rf_ram.memory\[27\]\[4\] _01516_ _01774_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08481__A1 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08207_ u_cpu.rf_ram.memory\[67\]\[5\] _03486_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09187_ u_cpu.rf_ram.memory\[127\]\[2\] _04120_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06399_ _02036_ _02038_ _02042_ _02044_ _01642_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08371__I _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08138_ _03415_ _03442_ _03447_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10040__A1 _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ _03337_ _03397_ _03402_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10100_ _04753_ _04782_ _04653_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11080_ _05468_ _05470_ _05472_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11889__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09733__A1 u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10031_ _02627_ _04699_ _04719_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08536__A2 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11540__A1 u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10343__A2 _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11982_ _00504_ net421 u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10933_ _05375_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _05335_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10297__B _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12603_ _01100_ net445 u_cpu.rf_ram.memory\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _03067_ _05158_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12514__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06066__I _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12534_ _01035_ net330 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05905__S0 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12465_ _00966_ net486 u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11359__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07098__S _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11416_ u_cpu.rf_ram.memory\[26\]\[5\] _05686_ _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08281__I _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12396_ _00897_ net474 u_cpu.rf_ram.memory\[115\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10031__A1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11347_ u_cpu.cpu.genblk3.csr.o_new_irq _05643_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08775__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__S0 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10582__A2 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ u_cpu.rf_ram.memory\[111\]\[1\] _05596_ _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _04889_ _04890_ _04893_ _04776_ _04695_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_13017_ _00078_ net532 u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11531__A1 _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10334__A2 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__I _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06669__C _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout282_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserv_2_542 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07440_ u_cpu.rf_ram.memory\[21\]\[4\] _02972_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07371_ _02902_ u_cpu.rf_ram_if.wdata0_r\[2\] _02917_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__12194__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09110_ u_cpu.rf_ram.memory\[12\]\[1\] _04066_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06322_ _01711_ _01968_ _01715_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08463__A1 u_cpu.rf_ram.memory\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10270__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ _04011_ _04016_ _04025_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06253_ _01552_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07018__A2 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06184_ _01576_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10226__I _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08766__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06321__S0 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09943_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _02726_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09715__A1 u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _04577_ _04578_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11522__A1 _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10325__A2 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08825_ _03888_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11057__I _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08756_ _03440_ _03183_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05968_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ _03137_ _03155_ _03158_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05899_ _01501_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08687_ _03746_ _03795_ _03802_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07638_ u_cpu.rf_ram.memory\[42\]\[3\] _03110_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06701__A1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _02940_ _03057_ _03064_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09308_ u_cpu.rf_ram.memory\[38\]\[4\] _04197_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _05144_ _05146_ u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08454__A1 u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12687__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10261__A1 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10261__B2 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09239_ _02905_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12250_ _00751_ net339 u_cpu.rf_ram.memory\[38\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07009__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08206__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11201_ u_cpu.rf_ram.memory\[10\]\[6\] _05543_ _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10013__A1 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09954__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12181_ _00695_ net374 u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06312__S0 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06768__A1 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11132_ _05475_ _05501_ _05506_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__A2 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11063_ u_cpu.rf_ram.memory\[107\]\[2\] _05461_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11513__A1 _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07445__I _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10014_ _04634_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06940__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11965_ _00487_ net28 u_cpu.rf_ram.memory\[53\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06379__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10916_ _05320_ _05363_ _05369_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08693__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11896_ _00418_ net270 u_cpu.rf_ram.memory\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10847_ u_cpu.rf_ram.memory\[28\]\[7\] _05311_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ u_cpu.rf_ram.memory\[95\]\[0\] _05284_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10252__A1 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12517_ _01018_ net307 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout128_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12448_ _00949_ net478 u_cpu.rf_ram.memory\[113\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10004__A1 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10046__I _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12379_ _00880_ net478 u_cpu.rf_ram.memory\[112\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06303__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06759__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout497_I net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06940_ _02517_ _02521_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06871_ _02486_ _02489_ _02494_ _02496_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06606__S1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05822_ _01440_ _01455_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08610_ _03754_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09590_ u_cpu.rf_ram.memory\[121\]\[3\] _04381_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08541_ _03661_ _03706_ _03708_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10866__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08472_ _03662_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11584__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07487__A2 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09881__B1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _02963_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10491__A1 _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06790__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07354_ _02876_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08436__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06305_ u_cpu.rf_ram.memory\[112\]\[2\] u_cpu.rf_ram.memory\[113\]\[2\] u_cpu.rf_ram.memory\[114\]\[2\]
+ u_cpu.rf_ram.memory\[115\]\[2\] _01679_ _01840_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08987__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _02763_ _02840_ _02841_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10794__A2 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _04014_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06236_ _01877_ _01879_ _01881_ _01883_ _01768_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06167_ u_cpu.rf_ram.memory\[52\]\[1\] u_cpu.rf_ram.memory\[53\]\[1\] u_cpu.rf_ram.memory\[54\]\[1\]
+ u_cpu.rf_ram.memory\[55\]\[1\] _01630_ _01631_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10546__A2 _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06098_ _01746_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ _04616_ _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09857_ _04566_ _04567_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ u_cpu.rf_ram.memory\[70\]\[1\] _03877_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06922__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _03283_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06773__I1 u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03730_ _03832_ _03834_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07478__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11750_ _00272_ net429 u_cpu.rf_ram.memory\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08096__I _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06525__I1 u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10701_ _04705_ _04974_ _04976_ _05227_ _04700_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10482__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11681_ _00203_ net389 u_cpu.rf_ram.memory\[51\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08427__A1 u_cpu.rf_ram.memory\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10632_ _04075_ _05172_ _05179_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10234__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _05136_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10234__B2 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06989__A1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10785__A2 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12302_ _00803_ net207 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ _03537_ _03083_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09927__A1 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12233_ _00008_ net285 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12164_ _00678_ net83 u_cpu.rf_ram.memory\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11115_ u_cpu.rf_ram.memory\[108\]\[4\] _05493_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12095_ _00609_ net336 u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11046_ u_cpu.rf_ram.memory\[106\]\[4\] _05448_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06764__I1 u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12852__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12997_ _00056_ net525 u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07469__A2 _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11948_ _00470_ net23 u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout245_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11879_ _00401_ net181 u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08418__A1 u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10225__A1 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout412_I net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10076__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08969__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09091__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ u_arbiter.i_wb_cpu_rdt\[19\] u_arbiter.i_wb_cpu_dbus_dat\[16\] _02671_ _02672_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12232__CLK net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06295__I3 u_cpu.rf_ram.memory\[111\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06021_ u_cpu.rf_ram.memory\[124\]\[0\] u_cpu.rf_ram.memory\[125\]\[0\] u_cpu.rf_ram.memory\[126\]\[0\]
+ u_cpu.rf_ram.memory\[127\]\[0\] _01668_ _01669_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09918__A1 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09394__A2 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12382__CLK net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07972_ _03329_ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06203__B _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09146__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06923_ _02492_ _02559_ _02560_ _02561_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout60_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09642_ _04413_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06854_ _02491_ _02493_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10700__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05805_ _01441_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06785_ _01604_ _02426_ _01640_ _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09573_ _04344_ _04365_ _04372_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11335__I _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06380__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08524_ _03693_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06429__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08455_ _03568_ _03650_ _03653_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06132__A2 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07406_ u_cpu.rf_ram_if.wdata1_r\[7\] _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08386_ u_cpu.rf_ram.memory\[60\]\[5\] _03601_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08409__A1 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07880__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10216__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07337_ _02885_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[2\] _02886_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09082__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06515__S0 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10767__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _02825_ _02818_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06164__I _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09007_ u_cpu.rf_ram.memory\[134\]\[3\] _04001_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06219_ _01540_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12725__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07199_ _02749_ u_scanchain_local.module_data_in\[51\] _02730_ u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout530 net532 net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_76_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12875__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _04600_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12920_ _01417_ net382 u_cpu.rf_ram.memory\[89\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08896__A1 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07723__I _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12851_ _01348_ net435 u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11802_ _00324_ net34 u_cpu.rf_ram.memory\[74\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12782_ _01279_ net112 u_cpu.rf_ram.memory\[84\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11733_ _00255_ net213 u_cpu.rf_ram.memory\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12255__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11664_ _00186_ net461 u_cpu.rf_ram.memory\[45\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07871__A2 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10207__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10615_ u_cpu.rf_ram.memory\[109\]\[6\] _05164_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09073__A1 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06506__S0 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11595_ _00117_ net212 u_cpu.rf_ram.memory\[81\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10758__A2 _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10546_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _05123_ _05125_ _02758_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08820__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07623__A2 _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10477_ _05081_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09376__A2 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12216_ _00730_ net343 u_cpu.rf_ram.memory\[125\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11183__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12147_ _00661_ net78 u_cpu.rf_ram.memory\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10930__A2 _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12078_ _00592_ net225 u_cpu.rf_ram.memory\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout195_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11029_ _05413_ _05433_ _05440_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10694__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout362_I net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__C _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06570_ u_cpu.rf_ram.memory\[12\]\[5\] u_cpu.rf_ram.memory\[13\]\[5\] u_cpu.rf_ram.memory\[14\]\[5\]
+ u_cpu.rf_ram.memory\[15\]\[5\] _01550_ _01553_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_79_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05960__I2 u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06693__B _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _03511_ _03496_ _03512_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ _02952_ _03458_ _03467_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11622__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10749__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ _02705_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08811__A1 u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07053_ u_arbiter.i_wb_cpu_rdt\[12\] u_arbiter.i_wb_cpu_dbus_dat\[9\] _02658_ _02662_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06004_ u_cpu.rf_ram.memory\[96\]\[0\] u_cpu.rf_ram.memory\[97\]\[0\] u_cpu.rf_ram.memory\[98\]\[0\]
+ u_cpu.rf_ram.memory\[99\]\[0\] _01652_ _01552_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07808__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11772__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07378__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11174__A2 _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07955_ u_cpu.rf_ram.memory\[17\]\[7\] _03313_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06906_ _02544_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08878__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07886_ _03274_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09625_ _04062_ _04402_ _04404_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06837_ _02473_ _02477_ u_arbiter.i_wb_cpu_dbus_we _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06353__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12278__CLK net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09556_ u_cpu.rf_ram.memory\[120\]\[6\] _04357_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06768_ _01692_ _02381_ _02390_ _02409_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_58_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08507_ u_cpu.rf_ram.memory\[56\]\[3\] _03686_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09487_ _04260_ _04310_ _04317_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06699_ _01580_ _02332_ _02341_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07302__A1 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05998__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08438_ _03640_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08374__I _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09055__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ u_cpu.rf_ram.memory\[61\]\[7\] _03583_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06108__B _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _05034_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11380_ u_cpu.cpu.genblk3.csr.o_new_irq _04242_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08802__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _04970_ _04983_ _04984_ _04985_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_106_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10262_ u_cpu.cpu.immdec.imm30_25\[5\] _04882_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07369__A1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12001_ _00006_ net292 u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10144__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _04695_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08030__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09933__I _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout360 net363 net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout371 net511 net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout382 net384 net382 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout393 net395 net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12903_ _01400_ net200 u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09530__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12834_ _01331_ net138 u_cpu.rf_ram.memory\[111\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12765_ _01262_ net171 u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08097__A2 _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__A1 u_cpu.rf_ram.memory\[123\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11716_ _00238_ net403 u_cpu.rf_ram.memory\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A2 _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12696_ _01193_ net153 u_cpu.rf_ram.memory\[102\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11647_ _00169_ net401 u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09046__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11795__CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11578_ _00100_ net213 u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout110_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10529_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _05116_ _05111_ _02725_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout208_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06670__I3 u_cpu.rf_ram.memory\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10054__I _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__A2 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09843__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06688__B _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07780__A1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07740_ u_cpu.rf_ram.memory\[51\]\[6\] _03174_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12420__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07671_ _03131_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09410_ _02899_ _03102_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06622_ _01971_ _02265_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06553_ _02187_ _02197_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09341_ u_cpu.rf_ram.memory\[36\]\[1\] _04218_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09285__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08088__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11092__A1 u_cpu.rf_ram.memory\[83\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08194__I _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06484_ u_cpu.rf_ram.memory\[36\]\[4\] u_cpu.rf_ram.memory\[37\]\[4\] u_cpu.rf_ram.memory\[38\]\[4\]
+ u_cpu.rf_ram.memory\[39\]\[4\] _01797_ _01680_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09272_ _04176_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07835__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _03494_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09037__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _03456_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09588__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11395__A2 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07105_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08085_ _03408_ _03410_ _03412_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08260__A2 _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07036_ u_arbiter.i_wb_cpu_rdt\[4\] _02651_ _02652_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06661__I3 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08012__A2 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08987_ u_cpu.rf_ram.memory\[135\]\[5\] _03986_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06574__A2 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07938_ _03313_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10658__A1 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07869_ u_cpu.rf_ram.memory\[4\]\[2\] _03263_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__I2 u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ u_cpu.rf_ram.memory\[8\]\[2\] _04393_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12913__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _05347_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05924__I2 u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09539_ _04350_ _04335_ _04351_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08079__A2 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__A1 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06709__S0 _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11083__A1 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12550_ _01050_ net173 u_cpu.rf_ram.memory\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11501_ _03646_ _05731_ _05740_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05837__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09028__A1 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12481_ _00982_ net240 u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11432_ u_cpu.rf_ram.memory\[25\]\[3\] _05698_ _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09579__A2 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11386__A2 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11363_ _05654_ u_cpu.cpu.genblk3.csr.mcause31 _05655_ _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08251__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07448__I _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06101__I2 u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _01439_ _04948_ _04968_ _04969_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11294_ _05606_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06652__I3 u_cpu.rf_ram.memory\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11138__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10245_ _04635_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08003__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12443__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10897__A1 u_cpu.rf_ram.memory\[101\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09751__A2 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _04788_ _04846_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__I3 u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06565__A2 _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__A1 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout190 net191 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07183__I _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10649__A1 u_cpu.rf_ram.memory\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A2 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07514__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11310__A2 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12593__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12817_ _01314_ net131 u_cpu.rf_ram.memory\[110\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout158_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11074__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12748_ _01245_ net115 u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05828__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout325_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12679_ _01176_ net47 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08490__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08742__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07358__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11129__A2 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08910_ _03754_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09890_ _04431_ _04585_ _04588_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07053__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09742__A2 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08841_ _03859_ _03890_ _03898_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06556__A2 _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07753__A1 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11810__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08772_ u_cpu.rf_ram.memory\[73\]\[4\] _03851_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05984_ _01629_ _01632_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07723_ _03167_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11301__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ _03018_ _03118_ _03121_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06605_ _01836_ _02248_ _01611_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09258__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ _03020_ _03070_ _03075_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11065__A1 u_cpu.rf_ram.memory\[107\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09324_ u_cpu.rf_ram.memory\[37\]\[2\] _04209_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06437__I _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06536_ u_cpu.rf_ram.memory\[72\]\[4\] u_cpu.rf_ram.memory\[73\]\[4\] u_cpu.rf_ram.memory\[74\]\[4\]
+ u_cpu.rf_ram.memory\[75\]\[4\] _01867_ _01695_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06167__S1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05819__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10812__A1 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _02925_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06467_ _01500_ _02111_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08481__A2 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _03420_ _03482_ _03489_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09186_ _04115_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06398_ _01926_ _02043_ _01929_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ u_cpu.rf_ram.memory\[75\]\[2\] _03446_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08233__A2 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09430__A1 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10040__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ u_cpu.rf_ram.memory\[77\]\[2\] _03401_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06795__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ _02611_ _02638_ _02639_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07044__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _04701_ _04712_ _04718_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09733__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06547__A2 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08099__I _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11981_ _00503_ net421 u_cpu.rf_ram.memory\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10932_ _05315_ _05376_ _05379_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10863_ _05338_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09249__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06570__I2 u_cpu.rf_ram.memory\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12602_ _01099_ net445 u_cpu.rf_ram.memory\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _05221_ _05284_ _05293_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06158__S1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12533_ _01034_ net329 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06791__B _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05905__S1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06483__A1 _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12464_ _00965_ net474 u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11415_ _05630_ _05682_ _05689_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12395_ _00896_ net481 u_cpu.rf_ram.memory\[115\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08224__A2 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07178__I _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06235__A1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06082__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11346_ u_cpu.cpu.decode.op21 _01442_ _01460_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06330__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11833__CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11277_ _05550_ _05595_ _05597_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13016_ _00077_ net532 u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09724__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _04891_ _04821_ _04892_ _04865_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07735__A1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _04831_ _04629_ _04732_ _04729_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11983__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout275_I net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_2_543 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08737__I _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A1 u_cpu.rf_ram.memory\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__S1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout442_I net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06710__A2 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11047__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ _02903_ u_cpu.rf_ram_if.wdata1_r\[2\] _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ u_cpu.rf_ram.memory\[84\]\[2\] u_cpu.rf_ram.memory\[85\]\[2\] u_cpu.rf_ram.memory\[86\]\[2\]
+ u_cpu.rf_ram.memory\[87\]\[2\] _01855_ _01713_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09660__A1 _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08463__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06252_ _01539_ _01898_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09040_ u_cpu.rf_ram.memory\[133\]\[7\] _04014_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12489__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _01660_ _01830_ _01663_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10558__B1 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06321__S1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07974__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09942_ _02705_ _04632_ _04633_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10443__S _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout90_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09715__A2 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09873_ u_arbiter.i_wb_cpu_rdt\[27\] _04495_ _04519_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11338__I _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11522__A2 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _03230_ _03887_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08755_ _03729_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05967_ _01514_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ u_cpu.rf_ram.memory\[44\]\[1\] _03156_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11286__A1 _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08686_ u_cpu.rf_ram.memory\[141\]\[4\] _03799_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05898_ _01512_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08151__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ _03020_ _03106_ _03111_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06701__A2 _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11038__A1 _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07568_ u_cpu.rf_ram.memory\[7\]\[5\] _03060_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11706__CLK net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04165_ _04193_ _04199_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06519_ u_cpu.rf_ram.memory\[116\]\[4\] u_cpu.rf_ram.memory\[117\]\[4\] u_cpu.rf_ram.memory\[118\]\[4\]
+ u_cpu.rf_ram.memory\[119\]\[4\] _02069_ _01685_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ _03014_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ _04101_ _04141_ _04150_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09403__A1 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ u_cpu.rf_ram.memory\[128\]\[3\] _04108_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08206__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11856__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11200_ _02978_ _05540_ _05547_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11210__A1 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10013__A2 _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12180_ _00694_ net192 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09954__A2 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07965__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__S1 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11131_ u_cpu.rf_ram.memory\[69\]\[2\] _05505_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09706__A2 _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11062_ _05456_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__A1 u_cpu.rf_ram.memory\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _04616_ _04690_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_23_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06940__A2 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11277__A1 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11964_ _00486_ net28 u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__A1 _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06379__S1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ u_cpu.rf_ram.memory\[102\]\[3\] _05367_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09890__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11895_ _00417_ net89 u_cpu.rf_ram.memory\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11029__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__I _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _05220_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10777_ _05282_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09388__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12516_ _01017_ net307 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12447_ _00948_ net481 u_cpu.rf_ram.memory\[113\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12781__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06059__I1 u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12378_ _00879_ net477 u_cpu.rf_ram.memory\[112\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07956__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06303__S1 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11329_ _02932_ _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12011__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout392_I net397 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06870_ _02497_ _02477_ _02503_ u_cpu.cpu.genblk3.csr.mstatus_mie _02509_ _02510_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08381__A1 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05821_ u_cpu.cpu.immdec.imm19_12_20\[8\] _01471_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11268__A1 _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08540_ u_cpu.rf_ram.memory\[54\]\[0\] _03707_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11729__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08471_ _03662_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09881__A1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08684__A2 _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06534__I2 u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07422_ _02871_ _02870_ _02893_ _02962_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_126_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__S1 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _02881_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08436__A2 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11879__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__I _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ _01836_ _01950_ _01676_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07284_ _02808_ u_scanchain_local.module_data_in\[66\] _02767_ u_arbiter.i_wb_cpu_dbus_adr\[29\]
+ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09023_ _04014_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06235_ _01763_ _01882_ _01756_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09936__A2 _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06166_ _01622_ _01813_ _01626_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06097_ _01745_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_105_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _04609_ _04611_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06470__I1 u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09856_ u_arbiter.i_wb_cpu_rdt\[21\] _04559_ _04560_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10703__B1 _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A1 _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06222__I1 u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _03843_ _03876_ _03878_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _02648_ _04512_ _04515_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06999_ _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06922__A2 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11259__A1 _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06773__I2 u_cpu.rf_ram.memory\[110\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08738_ u_cpu.rf_ram.memory\[72\]\[0\] _03833_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12654__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _03749_ _03784_ _03791_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10700_ _04645_ _04709_ _04732_ _04660_ _04974_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06686__A1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06230__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11680_ _00202_ net391 u_cpu.rf_ram.memory\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10482__A2 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10631_ u_cpu.rf_ram.memory\[3\]\[4\] _05176_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09624__A1 u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08427__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11431__A1 _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10234__A2 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10562_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _05130_ _05132_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12301_ _00802_ net197 u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06989__A2 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10493_ _05093_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12034__CLK net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12232_ _00020_ net281 u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06297__S0 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12163_ _00677_ net82 u_cpu.rf_ram.memory\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06360__I _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11114_ _05478_ _05489_ _05495_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12094_ _00608_ net337 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12184__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11498__A1 u_cpu.rf_ram.memory\[98\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ _05409_ _05444_ _05450_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09671__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10170__A1 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06913__A2 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12996_ _00055_ net525 u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11947_ _00469_ net23 u_cpu.rf_ram.memory\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__A2 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11878_ _00400_ net181 u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10829_ _05315_ _05312_ _05316_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09615__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout238_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11422__A1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09091__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout405_I net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__I _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06020_ _01618_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__A1 u_cpu.rf_ram.memory\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06288__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12527__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07366__I _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _03336_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__B _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09710_ _03012_ _04426_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06922_ u_cpu.cpu.alu.i_rs1 _02478_ _01452_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09581__I _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _03067_ _04179_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06853_ _02492_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05804_ _01447_ _01450_ _01454_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_3_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09572_ u_cpu.rf_ram.memory\[118\]\[4\] _04369_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06784_ u_cpu.rf_ram.memory\[116\]\[7\] u_cpu.rf_ram.memory\[117\]\[7\] u_cpu.rf_ram.memory\[118\]\[7\]
+ u_cpu.rf_ram.memory\[119\]\[7\] _02069_ _01638_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08523_ _03666_ _03694_ _03697_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08657__A2 _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06668__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__S0 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ u_cpu.rf_ram.memory\[58\]\[1\] _03651_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07405_ _02909_ _02946_ _02947_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08385_ _03575_ _03597_ _03604_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08409__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12057__CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11413__A1 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ u_cpu.rf_ram_if.rcnt\[0\] _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09082__A2 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06515__S1 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07093__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07267_ _02826_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _03742_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06218_ _01862_ _01864_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06840__A1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07198_ _02769_ _02765_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06149_ _01583_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout520 net523 net520 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout531 net532 net531 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _04599_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07148__A2 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09839_ _04553_ _04554_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10152__A1 _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06746__I2 u_cpu.rf_ram.memory\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12850_ _01347_ net436 u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11801_ _00323_ net34 u_cpu.rf_ram.memory\[74\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12781_ _01278_ net102 u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06659__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11732_ _00254_ net218 u_cpu.rf_ram.memory\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _00185_ net461 u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10614_ _04814_ _05161_ _05168_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06355__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11594_ _00116_ net212 u_cpu.rf_ram.memory\[81\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09073__A2 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06506__S1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10545_ _05126_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06131__I0 u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__A1 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10476_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[30\] _05078_
+ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12215_ _00729_ net343 u_cpu.rf_ram.memory\[125\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11574__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06304__B _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06434__I1 u_cpu.rf_ram.memory\[81\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12146_ _00660_ net82 u_cpu.rf_ram.memory\[133\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10391__A1 u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ _00591_ net222 u_cpu.rf_ram.memory\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06690__S0 _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11028_ u_cpu.rf_ram.memory\[105\]\[5\] _05436_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10143__A1 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout188_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__S0 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06898__A1 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10694__A2 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12979_ _00036_ net514 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05960__I3 u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__A2 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout522_I net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11171__I _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08170_ u_cpu.rf_ram.memory\[6\]\[7\] _03456_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05873__A2 _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07121_ u_cpu.cpu.genblk1.align.ctrl_misal _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08811__A2 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ _02661_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11917__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06003_ _01548_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10515__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10382__A1 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07954_ _03226_ _03315_ _03323_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06681__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06905_ _02468_ _02540_ _02543_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02544_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_56_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10134__A1 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07885_ _02726_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_95_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09624_ u_cpu.rf_ram.memory\[11\]\[0\] _04403_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06836_ u_cpu.rf_ram_if.rtrig1 _02475_ _02476_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__10685__A2 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09555_ _04346_ _04354_ _04361_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06767_ _01493_ _02399_ _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_55_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06884__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08506_ _03668_ _03682_ _03687_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ u_cpu.rf_ram.memory\[35\]\[5\] _04313_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08655__I _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06698_ _02334_ _02336_ _02338_ _02340_ _02072_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_19_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08437_ _02938_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11081__I _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ _03579_ _03585_ _03593_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09055__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07319_ _02484_ _01459_ _02869_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ _03509_ _03540_ _03548_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08802__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10330_ u_cpu.cpu.immdec.imm19_12_20\[5\] _04970_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06813__A1 _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12842__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ _04759_ _04918_ _04922_ _04698_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07369__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08566__A1 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12000_ _00005_ net292 u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10192_ _04843_ _04858_ _04859_ _04860_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10373__A1 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05963__B _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06672__S0 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12992__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout350 net352 net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08318__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout361 net363 net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06592__A3 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout372 net377 net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_98_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout383 net384 net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout394 net395 net394 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_12902_ _01399_ net195 u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06424__S0 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12222__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12833_ _01330_ net133 u_cpu.rf_ram.memory\[111\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06195__I3 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12764_ _01261_ net171 u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09294__A2 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11715_ _00237_ net403 u_cpu.rf_ram.memory\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12695_ _01192_ net153 u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06352__I0 u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06501__B1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11646_ _00168_ net401 u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11577_ _00099_ net209 u_cpu.rf_ram.memory\[82\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06804__A1 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10528_ _05107_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout103_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _05071_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06407__I1 u_cpu.rf_ram.memory\[109\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05873__B _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12129_ _00643_ net259 u_cpu.rf_ram.memory\[135\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06663__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08309__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07780__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout472_I net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10116__A1 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11166__I _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06415__S0 _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ _02957_ _03081_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06621_ u_cpu.rf_ram.memory\[64\]\[5\] u_cpu.rf_ram.memory\[65\]\[5\] u_cpu.rf_ram.memory\[66\]\[5\]
+ u_cpu.rf_ram.memory\[67\]\[5\] _01731_ _01972_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12715__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09340_ _04152_ _04217_ _04219_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06552_ _02190_ _02192_ _02194_ _02196_ _01768_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08475__I _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09285__A2 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ _02949_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06483_ _02121_ _02123_ _02125_ _02127_ _01578_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11092__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__I0 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06209__B _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ _03336_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout16_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12865__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08153_ _03456_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07104_ _02690_ _02643_ _02691_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08796__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ u_cpu.rf_ram.memory\[74\]\[0\] _03411_ _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07035_ _02633_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10245__I _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06654__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _03937_ _03982_ _03989_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07937_ _02964_ _02985_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10658__A2 _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07868_ _03258_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__A2 _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__I3 u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09607_ _04388_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06819_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_44_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12395__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ _03211_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ u_cpu.rf_ram.memory\[117\]\[7\] _04333_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09276__A2 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__S1 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09469_ _04262_ _04298_ _04306_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11083__A2 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11500_ u_cpu.rf_ram.memory\[98\]\[7\] _05729_ _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05837__A2 _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12480_ _00981_ net240 u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09028__A2 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11431_ _05625_ _05694_ _05699_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08787__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__B1 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11362_ _04228_ _02507_ _02515_ _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10594__A1 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10313_ u_cpu.cpu.immdec.imm19_12_20\[5\] _04670_ _04947_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06101__I3 u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13020__CLK net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11293_ _05512_ _03053_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10244_ _04904_ _04907_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06645__S0 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10175_ u_cpu.cpu.immdec.imm24_20\[1\] _04843_ _04844_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout180 net193 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11612__CLK net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout191 net192 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10649__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__A2 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08711__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06573__I0 u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12816_ _01313_ net132 u_cpu.rf_ram.memory\[110\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11762__CLK net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11074__A2 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12747_ _01244_ net116 u_cpu.rf_ram.memory\[106\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05828__A2 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12678_ _01175_ net50 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09019__A2 _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout220_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ _00151_ net209 u_cpu.rf_ram.memory\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout318_I net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06543__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07450__A1 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10337__A1 _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ u_cpu.rf_ram.memory\[143\]\[6\] _03893_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06636__S0 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07374__I _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _03745_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05983_ u_cpu.rf_ram.memory\[52\]\[0\] u_cpu.rf_ram.memory\[53\]\[0\] u_cpu.rf_ram.memory\[54\]\[0\]
+ u_cpu.rf_ram.memory\[55\]\[0\] _01630_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06211__C _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ _03084_ _02870_ _02962_ _03085_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_66_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ u_cpu.rf_ram.memory\[46\]\[1\] _03119_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06604_ u_cpu.rf_ram.memory\[120\]\[5\] u_cpu.rf_ram.memory\[121\]\[5\] u_cpu.rf_ram.memory\[122\]\[5\]
+ u_cpu.rf_ram.memory\[123\]\[5\] _01606_ _01837_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__B _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07584_ u_cpu.rf_ram.memory\[80\]\[2\] _03074_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09323_ _04204_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06535_ _01862_ _02179_ _01865_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05819__A2 _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09254_ _04161_ _04154_ _04163_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10812__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06466_ u_cpu.rf_ram.memory\[28\]\[4\] u_cpu.rf_ram.memory\[29\]\[4\] u_cpu.rf_ram.memory\[30\]\[4\]
+ u_cpu.rf_ram.memory\[31\]\[4\] _01504_ _01771_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08205_ u_cpu.rf_ram.memory\[67\]\[4\] _03486_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09185_ _04088_ _04116_ _04119_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06397_ u_cpu.rf_ram.memory\[48\]\[3\] u_cpu.rf_ram.memory\[49\]\[3\] u_cpu.rf_ram.memory\[50\]\[3\]
+ u_cpu.rf_ram.memory\[51\]\[3\] _01636_ _01927_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07549__I _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09965__S _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03441_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09430__A2 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07441__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08067_ _03396_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07018_ _02495_ _02629_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09194__A1 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11635__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07044__I1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__A1 u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08969_ u_cpu.rf_ram.memory\[136\]\[6\] _03974_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11980_ _00502_ net221 u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11785__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ u_cpu.rf_ram.memory\[103\]\[1\] _05377_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10500__A1 _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06555__I0 u_cpu.rf_ram.memory\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10862_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _05335_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12601_ _01098_ net446 u_cpu.rf_ram.memory\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06307__I0 u_cpu.rf_ram.memory\[116\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ u_cpu.rf_ram.memory\[95\]\[7\] _05282_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12532_ _01033_ net325 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10803__A2 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12463_ _00964_ net263 u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11414_ u_cpu.rf_ram.memory\[26\]\[4\] _05686_ _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12410__CLK net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12394_ _00895_ net491 u_cpu.rf_ram.memory\[115\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09421__A2 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11345_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06235__A2 _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11276_ u_cpu.rf_ram.memory\[111\]\[0\] _05596_ _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10319__A1 _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05994__B2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13015_ _00076_ net532 u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09185__A1 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06618__S0 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10227_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _04773_ _04892_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12560__CLK net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07194__I _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08932__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06389__I3 u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _04637_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _04759_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09488__A2 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout170_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserv_2_544 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__11444__I _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout268_I net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__B2 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11047__A2 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06561__I3 u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout435_I net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ _01852_ _01966_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07266__A4 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06251_ u_cpu.rf_ram.memory\[4\]\[2\] u_cpu.rf_ram.memory\[5\]\[2\] u_cpu.rf_ram.memory\[6\]\[2\]
+ u_cpu.rf_ram.memory\[7\]\[2\] _01782_ _01897_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06474__A2 _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12090__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06182_ u_cpu.rf_ram.memory\[104\]\[1\] u_cpu.rf_ram.memory\[105\]\[1\] u_cpu.rf_ram.memory\[106\]\[1\]
+ u_cpu.rf_ram.memory\[107\]\[1\] _01661_ _01571_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12903__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _04603_ u_arbiter.i_wb_cpu_rdt\[11\] _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09176__A1 _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09872_ u_arbiter.i_wb_cpu_dbus_dat\[27\] _04521_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout83_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09971__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _03369_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10730__A1 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08754_ _03755_ _03833_ _03842_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05966_ _01581_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07705_ _03129_ _03155_ _03157_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _03743_ _03795_ _03801_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05897_ _01539_ _01545_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08151__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07636_ u_cpu.rf_ram.memory\[42\]\[2\] _03110_ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07567_ _02934_ _03056_ _03063_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11038__A2 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09759__I _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09306_ u_cpu.rf_ram.memory\[38\]\[3\] _04197_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06518_ _02065_ _02162_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07498_ _03014_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12433__CLK net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09651__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ u_cpu.rf_ram.memory\[125\]\[7\] _04139_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07662__A1 u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06449_ _01735_ _02094_ _01738_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09168_ _04090_ _04104_ _04109_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09403__A2 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07414__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08119_ _03418_ _03429_ _03435_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11210__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12583__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ _04009_ _04052_ _04060_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06768__A3 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11130_ _05500_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09167__A1 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ _05404_ _05457_ _05460_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07717__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _04700_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08390__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ _00485_ net28 u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10914_ _05317_ _05363_ _05368_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11894_ _00416_ net89 u_cpu.rf_ram.memory\[61\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09890__A2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10845_ _05326_ _05313_ _05327_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11029__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10776_ _05282_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10788__A1 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06000__S1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07653__A1 u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12515_ _01016_ net307 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06700__I0 u_cpu.rf_ram.memory\[92\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11800__CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12446_ _00947_ net475 u_cpu.rf_ram.memory\[113\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07405__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11201__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__I2 u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12377_ _00878_ net477 u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07956__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11328_ _05628_ _05620_ _05629_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06821__I _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11950__CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09158__A1 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11259_ _05555_ _05583_ _05586_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__A1 u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout385_I net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10712__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12306__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ _01440_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08381__A2 _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11268__A2 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05990__I1 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09330__A1 u_cpu.rf_ram.memory\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06268__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08470_ _03550_ _03183_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12456__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09881__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07421_ _02895_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06534__I3 u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06695__A2 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10228__B1 _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07352_ _02900_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10779__A1 _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09633__A2 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05900__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06303_ u_cpu.rf_ram.memory\[120\]\[2\] u_cpu.rf_ram.memory\[121\]\[2\] u_cpu.rf_ram.memory\[122\]\[2\]
+ u_cpu.rf_ram.memory\[123\]\[2\] _01673_ _01837_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06447__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11440__A2 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10518__I _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _02837_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ _02961_ _04013_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06234_ u_cpu.rf_ram.memory\[140\]\[1\] u_cpu.rf_ram.memory\[141\]\[1\] u_cpu.rf_ram.memory\[142\]\[1\]
+ u_cpu.rf_ram.memory\[143\]\[1\] _01764_ _01765_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09397__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10454__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06165_ u_cpu.rf_ram.memory\[56\]\[1\] u_cpu.rf_ram.memory\[57\]\[1\] u_cpu.rf_ram.memory\[58\]\[1\]
+ u_cpu.rf_ram.memory\[59\]\[1\] _01623_ _01812_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07947__A2 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ _01514_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10951__A1 u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09149__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _04613_ _04615_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06470__I2 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09944__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09855_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _04557_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10703__A1 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10703__B2 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A2 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08806_ u_cpu.rf_ram.memory\[70\]\[0\] _03877_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06998_ _02621_ u_cpu.cpu.state.ibus_cyc _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09786_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _04507_ _04514_ _04486_ _04511_ _04515_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11259__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05949_ _01510_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08737_ _03831_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11084__I _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08668_ u_cpu.rf_ram.memory\[142\]\[5\] _03787_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09872__A2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07619_ u_cpu.rf_ram.memory\[78\]\[6\] _03093_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06230__S1 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10482__A3 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08599_ u_cpu.rf_ram.memory\[52\]\[4\] _03740_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10219__B1 _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12949__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10630_ _04073_ _05172_ _05178_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06906__I _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09624__A2 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05810__I u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _05135_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11431__A2 _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12300_ _00801_ net315 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10492_ _02635_ _05092_ _05089_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12231_ _00019_ net281 u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11195__A1 u_cpu.rf_ram.memory\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10242__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08060__A1 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12162_ _00676_ net85 u_cpu.rf_ram.memory\[131\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06297__S1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11113_ u_cpu.rf_ram.memory\[108\]\[3\] _05493_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12093_ _00607_ net336 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06461__I2 u_cpu.rf_ram.memory\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11044_ u_cpu.rf_ram.memory\[106\]\[3\] _05448_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11498__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__A2 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09560__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12479__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10170__A2 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12995_ _00054_ net521 u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10112__B _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11946_ _00468_ net37 u_cpu.rf_ram.memory\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07874__A1 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11877_ _00399_ net182 u_cpu.rf_ram.memory\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ u_cpu.rf_ram.memory\[28\]\[1\] _05313_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09615__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07626__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11422__A2 _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout133_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10759_ _05196_ _05271_ _05273_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09379__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout300_I net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12429_ _00930_ net49 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06288__S1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08051__A1 u_cpu.rf_ram.memory\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07970_ _02919_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06921_ _02485_ _02559_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09551__A1 _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _04081_ _04403_ _04412_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06852_ u_cpu.cpu.bne_or_bge _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08478__I _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07382__I _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05803_ _01453_ _01445_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_110_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09571_ _04342_ _04365_ _04371_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06783_ _02065_ _02424_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11846__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08106__A2 _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ u_cpu.rf_ram.memory\[55\]\[1\] _03695_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout46_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _03563_ _03650_ _03652_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07865__A1 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__S1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07404_ u_cpu.rf_ram.memory\[82\]\[6\] _02922_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08384_ u_cpu.rf_ram.memory\[60\]\[4\] _03601_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09102__I _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05971__S0 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07617__A1 u_cpu.rf_ram.memory\[78\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _02879_ _02883_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__11413__A2 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ _02824_ _02825_ _02819_ _02812_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_87_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09005_ _04000_ _03995_ _04002_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06217_ _01555_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07197_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11177__A1 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06148_ _01628_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08042__A1 u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10924__A1 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__A1 _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06079_ _01555_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout510 net511 net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09917__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout521 net523 net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_28_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout532 net536 net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09907_ _04598_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12621__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09838_ u_arbiter.i_wb_cpu_rdt\[16\] _04546_ _04547_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10152__A2 _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06746__I3 u_cpu.rf_ram.memory\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09769_ _02649_ _02651_ _04487_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11800_ _00322_ net34 u_cpu.rf_ram.memory\[74\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11101__A1 u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12780_ _01277_ net102 u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_92_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11731_ _00253_ net218 u_cpu.rf_ram.memory\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A1 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11662_ _00184_ net463 u_cpu.rf_ram.memory\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09012__I _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10613_ u_cpu.rf_ram.memory\[109\]\[5\] _05164_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10158__I _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11593_ _00115_ net410 u_cpu.rf_ram.memory\[81\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10207__A3 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10544_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _05123_ _05125_ u_cpu.cpu.ctrl.o_ibus_adr\[11\]
+ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12151__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__A2 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10475_ _05080_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11168__A1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11719__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12214_ _00728_ net299 u_cpu.rf_ram.memory\[125\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10915__A1 u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12145_ _00659_ net77 u_cpu.rf_ram.memory\[133\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10391__A2 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12076_ _00590_ net219 u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06690__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11869__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11027_ _05411_ _05432_ _05439_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09533__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11340__A1 _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10143__A2 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06737__I3 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__S1 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06898__A2 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05945__I1 u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12978_ _00035_ net514 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout250_I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11929_ _00451_ net74 u_cpu.rf_ram.memory\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout348_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05953__S0 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10068__I _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout515_I net518 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07120_ _02664_ _02703_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10454__I0 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08272__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08761__I _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07051_ u_arbiter.i_wb_cpu_rdt\[11\] u_arbiter.i_wb_cpu_dbus_dat\[8\] _02658_ _02661_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11159__A1 _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06002_ _01511_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__A1 u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ u_cpu.rf_ram.memory\[17\]\[6\] _03318_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06681__S1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09524__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08327__A2 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10531__I _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _02541_ _02542_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07884_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07326__B _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11331__A1 _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10134__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09623_ _04401_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06835_ u_cpu.rf_ram_if.rdata1\[0\] u_cpu.rf_ram_if.rtrig1 _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06766_ _02401_ _02403_ _02405_ _02407_ _01489_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09554_ u_cpu.rf_ram.memory\[120\]\[5\] _04357_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12024__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07840__I _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ u_cpu.rf_ram.memory\[56\]\[2\] _03686_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07838__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09485_ _04258_ _04309_ _04316_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06697_ _01604_ _02339_ _01640_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08436_ _03638_ _03624_ _03639_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ u_cpu.rf_ram.memory\[61\]\[6\] _03588_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07318_ _02618_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08298_ u_cpu.rf_ram.memory\[29\]\[6\] _03543_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10070__A1 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07249_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] u_cpu.cpu.ctrl.o_ibus_adr\[22\] u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _02802_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06813__A2 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06405__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _04920_ _04921_ _04824_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08015__A1 u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ u_cpu.cpu.immdec.imm24_20\[3\] _04843_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10373__A2 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06672__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout340 net341 net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08318__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout351 net352 net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout362 net363 net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout373 net377 net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout384 net385 net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06140__B _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout395 net397 net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12901_ _01398_ net437 u_cpu.rf_ram.memory\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06424__S1 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12832_ _01329_ net133 u_cpu.rf_ram.memory\[111\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12763_ _01260_ net186 u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12517__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11714_ _00236_ net462 u_cpu.rf_ram.memory\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12694_ _01191_ net153 u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06352__I1 u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06501__B2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11645_ _00167_ net164 u_cpu.rf_ram.memory\[78\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08581__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12667__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__A1 _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11576_ _00098_ net210 u_cpu.rf_ram.memory\[82\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10527_ _05115_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _05066_
+ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11691__CLK net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08557__A2 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06407__I2 u_cpu.rf_ram.memory\[110\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10389_ u_cpu.rf_ram.memory\[32\]\[6\] _05027_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11561__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10364__A2 _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06112__S0 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12128_ _00642_ net259 u_cpu.rf_ram.memory\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06663__S1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout298_I net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12059_ _00573_ net15 u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout465_I net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__S1 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _02257_ _02259_ _02261_ _02263_ _01858_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06551_ _01992_ _02195_ _01574_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12197__CLK net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10300__B _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09270_ _04174_ _04155_ _04175_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06482_ _01468_ _02126_ _01792_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08493__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06343__I1 u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08221_ _03498_ _03495_ _03499_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09587__I _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08152_ _03455_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08491__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08245__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07103_ _02630_ u_scanchain_local.module_data_in\[35\] _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10052__A1 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ _03409_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07034_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09745__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11552__A1 u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10355__A2 _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06654__S1 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ u_cpu.rf_ram.memory\[135\]\[4\] _03986_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07936_ _03228_ _03303_ _03312_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11304__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ _02915_ _03259_ _03262_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09606_ _04068_ _04389_ _04392_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06818_ _01476_ _02410_ _02459_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07798_ _02920_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _04176_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06749_ u_cpu.rf_ram.memory\[36\]\[7\] u_cpu.rf_ram.memory\[37\]\[7\] u_cpu.rf_ram.memory\[38\]\[7\]
+ u_cpu.rf_ram.memory\[39\]\[7\] _01679_ _01680_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09468_ u_cpu.rf_ram.memory\[92\]\[6\] _04301_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08419_ _03621_ _03624_ _03626_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__B2 _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09399_ u_cpu.rf_ram.memory\[91\]\[4\] _04254_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11430_ u_cpu.rf_ram.memory\[25\]\[2\] _05698_ _05699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10043__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__A1 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _01461_ _02512_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08787__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__B2 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10312_ _04664_ _04612_ _04967_ _04787_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11292_ _05568_ _05596_ _05605_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09736__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10243_ u_cpu.cpu.immdec.imm30_25\[3\] _04880_ _04905_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _04906_ _04683_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10346__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _04771_ _04845_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06645__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout170 net171 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06970__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout181 net184 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout192 net193 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11907__CLK net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__I1 u_cpu.rf_ram.memory\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12815_ _01312_ net131 u_cpu.rf_ram.memory\[110\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06096__I _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12746_ _01243_ net116 u_cpu.rf_ram.memory\[106\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A1 _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12677_ _01174_ net234 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11628_ _00150_ net217 u_cpu.rf_ram.memory\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08778__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout213_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11559_ _03643_ _05767_ _05775_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06789__A1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07450__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09727__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11534__A1 u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06636__S1 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08770_ _03853_ _03845_ _03854_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05982_ _01600_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06961__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07721_ _02884_ _03051_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06013__I0 u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08702__A2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07652_ _03010_ _03118_ _03120_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06564__I1 u_cpu.rf_ram.memory\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _01582_ _02246_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07583_ _03069_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07323__C _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04158_ _04205_ _04208_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06534_ u_cpu.rf_ram.memory\[68\]\[4\] u_cpu.rf_ram.memory\[69\]\[4\] u_cpu.rf_ram.memory\[70\]\[4\]
+ u_cpu.rf_ram.memory\[71\]\[4\] _01712_ _01863_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08466__A1 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10273__A1 _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06465_ _01497_ _02047_ _02110_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ u_cpu.rf_ram.memory\[124\]\[2\] _04162_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08204_ _03418_ _03482_ _03488_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08218__A1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09184_ u_cpu.rf_ram.memory\[127\]\[1\] _04117_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06396_ _02039_ _02041_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08769__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ _03413_ _03442_ _03445_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09430__A3 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ _03334_ _03397_ _03400_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07441__A2 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09718__A1 u_cpu.rf_ram.memory\[116\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07017_ _02492_ _02612_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11525__A1 u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09194__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06627__S1 _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10205__B _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08941__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _03939_ _03971_ _03978_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06952__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07919_ _03301_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08899_ u_cpu.rf_ram.memory\[39\]\[3\] _03933_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10930_ _05309_ _05376_ _05378_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10500__A2 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _05337_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12600_ _01097_ net446 u_cpu.rf_ram.memory\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08457__A1 u_cpu.rf_ram.memory\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10792_ _05218_ _05284_ _05292_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06307__I1 u_cpu.rf_ram.memory\[117\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10264__A1 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12531_ _01032_ net324 u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12462_ _00963_ net253 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11413_ _05628_ _05682_ _05688_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12393_ _00894_ net482 u_cpu.rf_ram.memory\[115\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06315__S0 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ _05640_ _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09709__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11275_ _05594_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11516__A1 u_cpu.rf_ram.memory\[100\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10319__A2 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05994__A2 _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13014_ _00075_ net531 u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09185__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _04645_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06618__S1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07196__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10157_ _04716_ _04641_ _04829_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06943__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ _02539_ _04699_ _04771_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_2_545 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout163_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__A2 _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08448__A1 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout330_I net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12729_ _01226_ net124 u_cpu.rf_ram.memory\[79\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout428_I net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__A1 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06250_ _01543_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09948__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06181_ _01656_ _01828_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09940_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11507__A1 u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09871_ _02683_ _04526_ _04576_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A1 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08923__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08822_ _03861_ _03877_ _03886_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout76_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08753_ u_cpu.rf_ram.memory\[72\]\[7\] _03831_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05965_ _01588_ _01597_ _01603_ _01612_ _01613_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_2_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07704_ u_cpu.rf_ram.memory\[44\]\[0\] _03156_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10869__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05896_ u_cpu.rf_ram.memory\[4\]\[0\] u_cpu.rf_ram.memory\[5\]\[0\] u_cpu.rf_ram.memory\[6\]\[0\]
+ u_cpu.rf_ram.memory\[7\]\[0\] _01542_ _01544_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08687__A1 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08684_ u_cpu.rf_ram.memory\[141\]\[3\] _03799_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10494__A1 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _03105_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13010__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08439__A1 u_cpu.rf_ram.memory\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07566_ u_cpu.rf_ram.memory\[7\]\[4\] _03060_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10246__A1 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09305_ _04161_ _04193_ _04198_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06517_ u_cpu.rf_ram.memory\[112\]\[4\] u_cpu.rf_ram.memory\[113\]\[4\] u_cpu.rf_ram.memory\[114\]\[4\]
+ u_cpu.rf_ram.memory\[115\]\[4\] _02066_ _01840_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07497_ _02964_ _03013_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09236_ _04099_ _04141_ _04149_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06448_ u_cpu.rf_ram.memory\[76\]\[3\] u_cpu.rf_ram.memory\[77\]\[3\] u_cpu.rf_ram.memory\[78\]\[3\]
+ u_cpu.rf_ram.memory\[79\]\[3\] _01979_ _01736_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_10_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06379_ u_cpu.rf_ram.memory\[32\]\[3\] u_cpu.rf_ram.memory\[33\]\[3\] u_cpu.rf_ram.memory\[34\]\[3\]
+ u_cpu.rf_ram.memory\[35\]\[3\] _01590_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09167_ u_cpu.rf_ram.memory\[128\]\[2\] _04108_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12728__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ u_cpu.rf_ram.memory\[76\]\[3\] _03433_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09098_ u_cpu.rf_ram.memory\[130\]\[6\] _04055_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08049_ u_cpu.rf_ram.memory\[139\]\[3\] _03388_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06413__B _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ u_cpu.rf_ram.memory\[107\]\[1\] _05458_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09167__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12878__CLK net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _04609_ _04653_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08678__A1 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11962_ _00484_ net37 u_cpu.rf_ram.memory\[54\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09015__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ u_cpu.rf_ram.memory\[102\]\[2\] _05367_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11893_ _00415_ net87 u_cpu.rf_ram.memory\[61\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06784__S0 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10844_ u_cpu.rf_ram.memory\[28\]\[6\] _05318_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12258__CLK net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _04295_ _03231_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06536__S0 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10788__A2 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12514_ _01015_ net307 u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A1 u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12445_ _00946_ net474 u_cpu.rf_ram.memory\[113\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__A2 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12376_ _00877_ net477 u_cpu.rf_ram.memory\[112\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ u_cpu.rf_ram.memory\[88\]\[3\] _05626_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09158__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ u_cpu.rf_ram.memory\[86\]\[1\] _05584_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10209_ _04874_ _04875_ _04861_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11189_ _02954_ _05539_ _05541_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06916__A1 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout378_I net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08669__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09330__A2 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ _02960_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08764__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07892__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__A1 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _02891_ _02899_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10228__B2 _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06527__S0 _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10779__A2 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06302_ _01667_ _01948_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07282_ _02836_ _02838_ _02839_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07644__A2 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06233_ _01758_ _01880_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09021_ _03369_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__A2 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11775__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06164_ _01592_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ _01691_ _01742_ _01743_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06080__A1 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09149__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _03274_ u_arbiter.i_wb_cpu_rdt\[15\] _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__I3 u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _04564_ _04565_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10703__A2 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _03875_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06222__I3 u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09785_ _04490_ _03283_ _04513_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06997_ net2 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08736_ _03831_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05948_ _01589_ _01594_ _01596_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12400__CLK net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08667_ _03746_ _03783_ _03790_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05879_ _01512_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ _03027_ _03090_ _03097_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08598_ _03745_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07549_ _03036_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10560_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _05130_ _05132_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08832__A1 u_cpu.rf_ram.memory\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _03131_ _03356_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _05084_ _05091_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12230_ _00018_ net287 u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07399__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11195__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10242__I1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12161_ _00675_ net79 u_cpu.rf_ram.memory\[131\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08060__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ _05475_ _05489_ _05494_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12092_ _00606_ net337 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06461__I3 u_cpu.rf_ram.memory\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11043_ _05406_ _05444_ _05449_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08899__A1 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09560__A2 _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A2 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A1 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12994_ _00053_ net521 u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11945_ _00467_ net37 u_cpu.rf_ram.memory\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11648__CLK net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07323__A1 _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08584__I _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07874__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11876_ _00398_ net181 u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10827_ _05201_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10758_ u_cpu.rf_ram.memory\[94\]\[0\] _05272_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10630__A1 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout126_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10689_ u_cpu.rf_ram.memory\[93\]\[6\] _05206_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12428_ _00929_ net47 u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12359_ _00860_ net441 u_cpu.rf_ram.memory\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08051__A2 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout495_I net509 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06920_ u_cpu.cpu.alu.i_rs1 _02478_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06851_ _02490_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09551__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10303__B _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05802_ _01451_ u_cpu.cpu.bne_or_bge _01452_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06279__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09570_ u_cpu.rf_ram.memory\[118\]\[3\] _04369_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06782_ u_cpu.rf_ram.memory\[112\]\[7\] u_cpu.rf_ram.memory\[113\]\[7\] u_cpu.rf_ram.memory\[114\]\[7\]
+ u_cpu.rf_ram.memory\[115\]\[7\] _02066_ _01631_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08521_ _03661_ _03694_ _03696_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12573__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08452_ u_cpu.rf_ram.memory\[58\]\[0\] _03651_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07865__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05911__I _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout39_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _02945_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09067__A1 u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08383_ _03573_ _03597_ _03603_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__S1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07334_ _02484_ _02880_ _02882_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07617__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__A1 _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__I0 u_cpu.rf_ram.memory\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10465__S _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09004_ u_cpu.rf_ram.memory\[134\]\[2\] _04001_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06216_ u_cpu.rf_ram.memory\[68\]\[1\] u_cpu.rf_ram.memory\[69\]\[1\] u_cpu.rf_ram.memory\[70\]\[1\]
+ u_cpu.rf_ram.memory\[71\]\[1\] _01725_ _01863_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07196_ _02763_ _02764_ _02765_ _02768_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_69_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__A2 _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06147_ _01493_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08042__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ u_cpu.rf_ram.memory\[68\]\[0\] u_cpu.rf_ram.memory\[69\]\[0\] u_cpu.rf_ram.memory\[70\]\[0\]
+ u_cpu.rf_ram.memory\[71\]\[0\] _01725_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout500 net501 net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__B u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout511 net512 net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09906_ _02632_ _02702_ _04597_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xfanout522 net523 net522 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout533 net536 net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_58_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09837_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _04544_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06356__A2 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12916__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06189__I _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _04490_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _03621_ _03820_ _03822_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09699_ _04433_ _04447_ _04452_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A2 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _00252_ net219 u_cpu.rf_ram.memory\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07856__A2 _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11661_ _00183_ net401 u_cpu.rf_ram.memory\[46\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10612_ _04812_ _05160_ _05167_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11592_ _00114_ net212 u_cpu.rf_ram.memory\[81\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06667__I0 u_cpu.rf_ram.memory\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10612__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _05110_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10463__I1 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10474_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _05078_
+ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11168__A2 _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12213_ _00727_ net298 u_cpu.rf_ram.memory\[125\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09230__A1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08033__A2 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12446__CLK net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07241__B1 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12144_ _00658_ net62 u_cpu.rf_ram.memory\[133\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12075_ _00589_ net222 u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11026_ u_cpu.rf_ram.memory\[105\]\[4\] _05436_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09533__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07544__A1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11340__A2 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12596__CLK net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06099__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12977_ _00034_ net516 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11928_ _00450_ net73 u_cpu.rf_ram.memory\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11859_ _00381_ net108 u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout243_I net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05953__S1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06658__I0 u_cpu.rf_ram.memory\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10603__A1 _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout410_I net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout508_I net509 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08272__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ _02660_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06001_ _01646_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11159__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__A2 _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__B1 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07083__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11813__CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07952_ _03224_ _03315_ _03322_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06511__B _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05906__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06903_ u_cpu.cpu.decode.opcode\[1\] _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09524__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07883_ _03271_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07535__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09622_ _04401_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06834_ u_cpu.rf_ram.rdata\[0\] _02474_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09553_ _04344_ _04353_ _04360_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06765_ _01698_ _02406_ _01654_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08504_ _03681_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09484_ u_cpu.rf_ram.memory\[35\]\[4\] _04313_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07838__A2 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06696_ u_cpu.rf_ram.memory\[116\]\[6\] u_cpu.rf_ram.memory\[117\]\[6\] u_cpu.rf_ram.memory\[118\]\[6\]
+ u_cpu.rf_ram.memory\[119\]\[6\] _02069_ _01638_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05849__A1 _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ u_cpu.rf_ram.memory\[5\]\[4\] _03632_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10842__A1 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ _03577_ _03585_ _03592_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06649__I0 u_cpu.rf_ram.memory\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11398__A2 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07317_ _02866_ _02868_ _02865_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09460__A1 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _03507_ _03540_ _03547_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06274__A1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12469__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09212__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07179_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _02745_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _02754_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09783__I _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07074__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ u_cpu.cpu.immdec.imm24_20\[4\] _04787_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout330 net331 net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05816__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout341 net342 net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout352 net353 net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout363 net367 net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout374 net376 net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XANTENNA__06329__A2 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout385 net386 net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12900_ _01397_ net437 u_cpu.rf_ram.memory\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout396 net397 net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12831_ _01328_ net132 u_cpu.rf_ram.memory\[111\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A1 u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11086__A1 u_cpu.rf_ram.memory\[83\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12762_ _01259_ net207 u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07829__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09023__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10833__A1 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11713_ _00235_ net462 u_cpu.rf_ram.memory\[47\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12693_ _01190_ net134 u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06501__A2 _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11644_ _00166_ net163 u_cpu.rf_ram.memory\[78\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10436__I1 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11575_ _00097_ net209 u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08254__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06265__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10526_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _05108_ _05111_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10118__B _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11836__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10457_ _05070_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09203__A1 _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08006__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07065__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _04814_ _05024_ _05031_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07765__A1 u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06112__S1 _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11561__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10364__A3 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12127_ _00641_ net258 u_cpu.rf_ram.memory\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09506__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12058_ _00572_ net16 u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08102__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout193_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07517__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05791__A3 u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11009_ _05413_ _05421_ _05428_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout360_I net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11463__I _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout458_I net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06550_ u_cpu.rf_ram.memory\[132\]\[4\] u_cpu.rf_ram.memory\[133\]\[4\] u_cpu.rf_ram.memory\[134\]\[4\]
+ u_cpu.rf_ram.memory\[135\]\[4\] _01993_ _02106_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ u_cpu.rf_ram.memory\[12\]\[4\] u_cpu.rf_ram.memory\[13\]\[4\] u_cpu.rf_ram.memory\[14\]\[4\]
+ u_cpu.rf_ram.memory\[15\]\[4\] _01550_ _01572_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09690__A1 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08493__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08220_ u_cpu.rf_ram.memory\[66\]\[1\] _03496_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08151_ _03050_ _03454_ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08245__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10588__B1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07388__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07102_ u_arbiter.i_wb_cpu_dbus_dat\[30\] _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ _03409_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07033_ _02648_ _02634_ _02650_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12761__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09745__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__A1 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11552__A2 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _03935_ _03982_ _03988_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07935_ u_cpu.rf_ram.memory\[16\]\[7\] _03301_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07508__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11304__A2 _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07866_ u_cpu.rf_ram.memory\[4\]\[1\] _03260_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08181__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09605_ u_cpu.rf_ram.memory\[8\]\[1\] _04390_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06817_ _02449_ _02458_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07797_ _03215_ _03212_ _03216_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12141__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11068__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09536_ _04348_ _04335_ _04349_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06748_ _02383_ _02385_ _02387_ _02389_ _01740_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_77_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11709__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10815__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09467_ _04260_ _04298_ _04305_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06679_ _01493_ _02312_ _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08484__A2 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08418_ u_cpu.rf_ram.memory\[5\]\[0\] _03625_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12291__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _04167_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ u_cpu.rf_ram.memory\[62\]\[7\] _03564_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08236__A2 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A2 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__A2 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _05650_ _05641_ _05653_ _02512_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07995__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _04740_ _04960_ _04961_ _04966_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_11291_ u_cpu.rf_ram.memory\[111\]\[7\] _05594_ _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07047__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09736__A2 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ u_arbiter.i_wb_cpu_rdt\[28\] u_arbiter.i_wb_cpu_rdt\[12\] _02709_ _04906_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ u_cpu.cpu.immdec.imm24_20\[0\] _04843_ _04844_ u_cpu.cpu.immdec.imm24_20\[1\]
+ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__I _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout160 net161 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout171 net179 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06970__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout182 net184 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout193 net230 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08172__A1 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11059__A1 _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12814_ _01311_ net131 u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12634__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10806__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12745_ _01242_ net115 u_cpu.rf_ram.memory\[106\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12676_ _01173_ net48 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _00149_ net217 u_cpu.rf_ram.memory\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08227__A2 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11558_ u_cpu.rf_ram.memory\[23\]\[6\] _05770_ _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09975__A2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06789__A2 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07986__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06333__S1 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ _04814_ _05096_ _05103_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout206_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11489_ _05729_ _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07038__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12014__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09727__A2 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07738__A1 u_cpu.rf_ram.memory\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11534__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05981_ _01583_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12164__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A2 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07720_ _03150_ _03156_ _03165_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07671__I _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08163__A1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ u_cpu.rf_ram.memory\[46\]\[0\] _03119_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06602_ u_cpu.rf_ram.memory\[124\]\[5\] u_cpu.rf_ram.memory\[125\]\[5\] u_cpu.rf_ram.memory\[126\]\[5\]
+ u_cpu.rf_ram.memory\[127\]\[5\] _01947_ _01707_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06287__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07582_ _03018_ _03070_ _03073_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ u_cpu.rf_ram.memory\[37\]\[1\] _04206_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06533_ _01971_ _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09663__A1 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10273__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout21_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06021__S0 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _04153_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06464_ _02098_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08203_ u_cpu.rf_ram.memory\[67\]\[3\] _03486_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08218__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ _04083_ _04116_ _04118_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06395_ u_cpu.rf_ram.memory\[52\]\[3\] u_cpu.rf_ram.memory\[53\]\[3\] u_cpu.rf_ram.memory\[54\]\[3\]
+ u_cpu.rf_ram.memory\[55\]\[3\] _01630_ _02040_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06229__A1 _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ u_cpu.rf_ram.memory\[75\]\[1\] _03443_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08065_ u_cpu.rf_ram.memory\[77\]\[1\] _03398_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07846__I _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07016_ _02637_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09718__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07729__A1 u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12507__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06088__S0 _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08967_ u_cpu.rf_ram.memory\[136\]\[5\] _03974_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06952__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07918_ _03301_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08898_ _03742_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12657__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07849_ u_cpu.rf_ram.memory\[50\]\[3\] _03249_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10860_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _05335_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ u_cpu.rf_ram.memory\[117\]\[1\] _04335_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10791_ u_cpu.rf_ram.memory\[95\]\[6\] _05287_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08457__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09654__A1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06307__I2 u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12530_ _01031_ net324 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11461__A1 _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10264__A2 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12461_ _00962_ net253 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09406__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08209__A2 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11412_ u_cpu.rf_ram.memory\[26\]\[3\] _05686_ _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11213__A1 _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12037__CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09957__A2 _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12392_ _00893_ net481 u_cpu.rf_ram.memory\[115\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06315__S1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11343_ _05638_ _05639_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09709__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11274_ _05594_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12187__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11516__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13013_ _00074_ net530 u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10225_ _04672_ _04781_ _04684_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10156_ _04764_ _04641_ _04709_ _04733_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__A2 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10087_ _04759_ _04760_ _04770_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_59_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09893__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xserv_2_546 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__A1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout156_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10989_ u_cpu.rf_ram.memory\[99\]\[6\] _05407_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06459__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12728_ _01225_ net128 u_cpu.rf_ram.memory\[79\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07120__A2 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12659_ _01156_ net236 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout323_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11204__A1 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__A2 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06180_ u_cpu.rf_ram.memory\[108\]\[1\] u_cpu.rf_ram.memory\[109\]\[1\] u_cpu.rf_ram.memory\[110\]\[1\]
+ u_cpu.rf_ram.memory\[111\]\[1\] _01549_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09948__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09870_ u_arbiter.i_wb_cpu_rdt\[26\] _04492_ _04574_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A2 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ u_cpu.rf_ram.memory\[70\]\[7\] _03875_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10820__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08752_ _03752_ _03833_ _03841_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05964_ _01576_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05914__I _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07703_ _03154_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _03739_ _03795_ _03800_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05895_ _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09884__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08687__A2 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07634_ _03018_ _03106_ _03109_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10494__A2 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07565_ _02928_ _03056_ _03062_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08439__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09636__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09304_ u_cpu.rf_ram.memory\[38\]\[2\] _04197_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06516_ _01836_ _02160_ _01611_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10246__A2 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ _03012_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07111__A2 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ u_cpu.rf_ram.memory\[125\]\[6\] _04144_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06447_ _01730_ _02092_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09939__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06870__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09166_ _04103_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ _01592_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06870__B2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ _03415_ _03429_ _03434_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _04007_ _04052_ _04059_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ _03337_ _03384_ _03389_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__I _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08375__A1 u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10010_ _04698_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09999_ _04650_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10182__A1 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06925__A2 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__S0 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08127__A1 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08200__I _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11961_ _00483_ net24 u_cpu.rf_ram.memory\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08678__A2 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10912_ _05362_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11892_ _00414_ net87 u_cpu.rf_ram.memory\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06784__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10843_ _05217_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09627__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10774_ _05221_ _05272_ _05281_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12513_ _01014_ net307 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06536__S1 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06700__I2 u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12444_ _00945_ net249 u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12375_ _00876_ net477 u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11577__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11326_ _02926_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06613__A1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06323__C _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11257_ _05550_ _05583_ _05585_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A1 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10208_ _04724_ _04686_ _04623_ _04688_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11188_ u_cpu.rf_ram.memory\[10\]\[0\] _05540_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10173__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10640__I _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ u_cpu.rf_ram.memory\[114\]\[5\] _04808_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12972__CLK net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08110__I _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout273_I net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__A2 _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12202__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07341__A2 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06775__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout440_I net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__A1 u_cpu.rf_ram.memory\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout538_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07350_ _02898_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10228__A2 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09094__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06527__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06301_ u_cpu.rf_ram.memory\[124\]\[2\] u_cpu.rf_ram.memory\[125\]\[2\] u_cpu.rf_ram.memory\[126\]\[2\]
+ u_cpu.rf_ram.memory\[127\]\[2\] _01947_ _01669_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06152__I0 u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07281_ _02808_ u_scanchain_local.module_data_in\[65\] _02767_ u_arbiter.i_wb_cpu_dbus_adr\[28\]
+ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12352__CLK net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _04011_ _03996_ _04012_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06232_ u_cpu.rf_ram.memory\[136\]\[1\] u_cpu.rf_ram.memory\[137\]\[1\] u_cpu.rf_ram.memory\[138\]\[1\]
+ u_cpu.rf_ram.memory\[139\]\[1\] _01759_ _01760_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08780__I _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _01615_ _01810_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07396__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05909__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06094_ _01475_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06080__A2 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09922_ _04603_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08357__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09853_ u_arbiter.i_wb_cpu_rdt\[20\] _04559_ _04560_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10164__A1 _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10164__B2 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _03875_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09784_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _04487_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06996_ _02614_ _02617_ _02619_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_58_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09116__I _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A2 _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ _03440_ _03328_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05947_ _01595_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08666_ u_cpu.rf_ram.memory\[142\]\[4\] _03787_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05878_ _01523_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07617_ u_cpu.rf_ram.memory\[78\]\[5\] _03093_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09609__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08597_ _02931_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ _02952_ _03040_ _03049_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09085__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06143__I0 u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07479_ _02969_ _02999_ _03002_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08832__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09218_ _04101_ _04129_ _04138_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06843__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _02874_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12845__CLK net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09149_ _04095_ _04085_ _04096_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08596__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12160_ _00674_ net84 u_cpu.rf_ram.memory\[131\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11111_ u_cpu.rf_ram.memory\[108\]\[2\] _05493_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12995__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12091_ _00605_ net337 u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11042_ u_cpu.rf_ram.memory\[106\]\[2\] _05448_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10155__A1 _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07020__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10460__I _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12225__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12993_ _00052_ net521 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11944_ _00466_ net67 u_cpu.rf_ram.memory\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11875_ _00397_ net181 u_cpu.rf_ram.memory\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10826_ _05309_ _05312_ _05314_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09076__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10757_ _05270_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07626__A3 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10630__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__I1 u_cpu.rf_ram.memory\[109\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10688_ _05217_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12427_ _00928_ net47 u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout119_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12358_ _00859_ net423 u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08105__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ u_cpu.rf_ram.memory\[87\]\[6\] _05611_ _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12289_ _00790_ net380 u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout390_I net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10146__A1 _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09000__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout488_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06850_ _01451_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10697__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10303__C _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ u_cpu.cpu.csr_d_sel _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_62_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ _01660_ _02422_ _01611_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08520_ u_cpu.rf_ram.memory\[55\]\[0\] _03695_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07314__A2 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08451_ _03649_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07402_ _02944_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ u_cpu.rf_ram.memory\[60\]\[3\] _03601_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11742__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09067__A2 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12868__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07333_ u_cpu.cpu.immdec.imm11_7\[1\] _02881_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08814__A2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06825__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07264_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06676__I1 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ _03994_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06215_ _01562_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07195_ _02766_ u_scanchain_local.module_data_in\[50\] _02767_ u_arbiter.i_wb_cpu_dbus_adr\[13\]
+ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06146_ _01784_ _01788_ _01790_ _01793_ _01578_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10385__A1 u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__A1 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ _01562_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout501 net503 net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12248__CLK net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09905_ _04596_ _02699_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout512 net5 net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10137__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout523 net524 net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout534 net535 net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_28_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07002__A1 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _04551_ _04552_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07553__A2 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _04489_ _04493_ _04498_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06979_ _02599_ _02593_ _02605_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ u_cpu.rf_ram.memory\[13\]\[0\] _03821_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ u_cpu.rf_ram.memory\[115\]\[2\] _04451_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08649_ _03641_ _03772_ _03779_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11660_ _00182_ net405 u_cpu.rf_ram.memory\[46\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09058__A2 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ u_cpu.rf_ram.memory\[109\]\[4\] _05164_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11591_ _00113_ net189 u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06667__I1 u_cpu.rf_ram.memory\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10542_ _05124_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10612__A2 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06131__I3 u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13023__CLK net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _05079_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12212_ _00726_ net294 u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09230__A2 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07241__A1 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12143_ _00657_ net44 u_cpu.rf_ram.memory\[133\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07241__B2 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12074_ _00588_ net67 u_cpu.rf_ram.memory\[143\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06601__C _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _05409_ _05432_ _05438_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12976_ _00033_ net514 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _00449_ net86 u_cpu.rf_ram.memory\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11858_ _00380_ net106 u_cpu.rf_ram.memory\[65\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10809_ u_cpu.rf_ram.memory\[96\]\[5\] _05299_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11789_ _00311_ net165 u_cpu.rf_ram.memory\[77\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout236_I net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10064__B1 _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10603__A2 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05887__C _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout403_I net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06283__A2 _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ u_cpu.rf_ram.memory\[100\]\[0\] u_cpu.rf_ram.memory\[101\]\[0\] u_cpu.rf_ram.memory\[102\]\[0\]
+ u_cpu.rf_ram.memory\[103\]\[0\] _01647_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10367__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07232__A1 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__A2 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07951_ u_cpu.rf_ram.memory\[17\]\[5\] _03318_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05794__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06902_ _02521_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12540__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07882_ _03270_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08732__A1 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07535__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09621_ _04400_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06833_ u_cpu.rf_ram.regzero _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_110_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09552_ u_cpu.rf_ram.memory\[120\]\[4\] _04357_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06764_ u_cpu.rf_ram.memory\[48\]\[7\] u_cpu.rf_ram.memory\[49\]\[7\] u_cpu.rf_ram.memory\[50\]\[7\]
+ u_cpu.rf_ram.memory\[51\]\[7\] _01699_ _01700_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05922__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _03666_ _03682_ _03685_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07299__A1 _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11095__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04256_ _04309_ _04315_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06695_ _02065_ _02337_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08434_ _03637_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05849__A2 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ u_cpu.rf_ram.memory\[61\]\[5\] _03588_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10476__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ _02867_ _02576_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06649__I1 u_cpu.rf_ram.memory\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08296_ u_cpu.rf_ram.memory\[29\]\[5\] _03543_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _02800_ _02802_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06274__A2 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12070__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _02752_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10358__A1 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09212__A2 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11638__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06129_ u_cpu.rf_ram.memory\[20\]\[1\] u_cpu.rf_ram.memory\[21\]\[1\] u_cpu.rf_ram.memory\[22\]\[1\]
+ u_cpu.rf_ram.memory\[23\]\[1\] _01524_ _01525_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07774__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__A1 u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout320 net321 net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout331 net332 net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout342 net354 net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout353 net354 net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout364 net366 net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11788__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout375 net377 net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07526__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout386 net409 net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _04531_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout397 net408 net397 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12830_ _01327_ net132 u_cpu.rf_ram.memory\[111\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11086__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12761_ _01258_ net207 u_cpu.rf_ram.memory\[83\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07252__C _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _00234_ net404 u_cpu.rf_ram.memory\[47\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12692_ _01189_ net136 u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11643_ _00165_ net164 u_cpu.rf_ram.memory\[78\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11574_ _00096_ net209 u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12413__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10597__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07462__A1 _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06265__A2 _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _05114_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _05066_
+ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10349__A1 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09203__A2 _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12563__CLK net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10387_ u_cpu.rf_ram.memory\[32\]\[5\] _05027_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12126_ _00640_ net258 u_cpu.rf_ram.memory\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08962__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12057_ _00571_ net9 u_cpu.rf_ram.memory\[71\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08714__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07517__A2 _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ u_cpu.rf_ram.memory\[79\]\[5\] _05424_ _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout186_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08190__A2 _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout353_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12959_ u_scanchain_local.module_data_in\[69\] net534 u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06480_ _01547_ _02124_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__B1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09690__A2 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout520_I net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07669__I _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08150_ _03453_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09442__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ _02689_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06256__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07453__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _03395_ _03102_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12906__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07032_ _02649_ _02609_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout99_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08953__A1 _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06803__I1 u_cpu.rf_ram.memory\[77\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08983_ u_cpu.rf_ram.memory\[135\]\[3\] _03986_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07934_ _03226_ _03303_ _03311_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__A2 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08705__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07865_ _02908_ _03259_ _03261_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09604_ _04062_ _04389_ _04391_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08181__A2 _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06816_ _02451_ _02453_ _02455_ _02457_ _01470_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07796_ u_cpu.rf_ram.memory\[48\]\[1\] _03213_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06747_ _01468_ _02388_ _01521_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11068__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09535_ u_cpu.rf_ram.memory\[117\]\[6\] _04340_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06582__I3 u_cpu.rf_ram.memory\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09130__A1 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ u_cpu.rf_ram.memory\[92\]\[5\] _04301_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06678_ _02314_ _02316_ _02318_ _02320_ _01489_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07141__B1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08417_ _03623_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07692__A1 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09397_ _04256_ _04248_ _04257_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ _03352_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09433__A2 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07444__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ u_cpu.rf_ram.memory\[64\]\[7\] _03525_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12586__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10310_ _04963_ _04965_ _04835_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11290_ _05566_ _05596_ _05604_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10241_ _04717_ _04879_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07047__I1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__A2 _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08944__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10172_ _04676_ _04841_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout150 net161 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout161 net162 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout172 net178 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout183 net184 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout194 net202 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10503__A1 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08172__A2 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06183__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11059__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12813_ _01310_ net131 u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06573__I3 u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09121__A1 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10806__A2 _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12744_ _01241_ net143 u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__A1 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12675_ _01172_ net48 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11803__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12929__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06393__I _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11626_ _00148_ net217 u_cpu.rf_ram.memory\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A1 _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06238__A2 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11231__A2 _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _03640_ _05767_ _05774_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07986__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ u_cpu.rf_ram.memory\[30\]\[5\] _05099_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11488_ _03627_ _05730_ _05733_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11953__CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10990__A1 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__A1 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout101_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07038__I1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10439_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _05060_
+ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07199__B1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06342__B _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12309__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12109_ _00623_ net293 u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05980_ _01628_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11298__A2 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout470_I net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08163__A2 _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09360__A1 _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _03117_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__I2 u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12459__CLK net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06601_ _02238_ _02240_ _02242_ _02244_ _01832_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_81_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07581_ u_cpu.rf_ram.memory\[80\]\[1\] _03071_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09320_ _04152_ _04205_ _04207_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06532_ u_cpu.rf_ram.memory\[64\]\[4\] u_cpu.rf_ram.memory\[65\]\[4\] u_cpu.rf_ram.memory\[66\]\[4\]
+ u_cpu.rf_ram.memory\[67\]\[4\] _01731_ _01972_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A2 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09251_ _04160_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06463_ _02100_ _02103_ _02105_ _02108_ _01768_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06021__S1 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11470__A2 _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08202_ _03415_ _03482_ _03487_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09182_ u_cpu.rf_ram.memory\[127\]\[0\] _04117_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout14_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06394_ _01600_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09415__A2 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _03408_ _03442_ _03444_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11222__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07977__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ _03326_ _03397_ _03399_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10981__A1 _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ _02632_ _02634_ _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09179__A1 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09119__I _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08926__A1 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06088__S1 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__I0 u_cpu.rf_ram.memory\[92\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10733__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ _03937_ _03970_ _03977_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07917_ _02964_ _03068_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11384__I _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08897_ _03932_ _03927_ _03934_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09351__A1 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07848_ _03217_ _03245_ _03250_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07779_ u_cpu.rf_ram.memory\[43\]\[3\] _03203_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09103__A1 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _04157_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10790_ _05215_ _05284_ _05291_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__A2 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__A1 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11461__A2 _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ u_cpu.cpu.state.init_done _04242_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12460_ _00961_ net253 u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__A2 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06146__C _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11411_ _05625_ _05682_ _05687_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07417__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12391_ _00892_ net481 u_cpu.rf_ram.memory\[115\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11213__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11342_ _02462_ _02507_ _02501_ _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11273_ _03230_ _05455_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07258__B _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09029__I _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08917__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10224_ _04644_ _04731_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09965__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13012_ _00073_ net530 u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10724__A1 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07196__A3 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ _04823_ _04827_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06943__A3 _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10086_ _04761_ _04769_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11294__I _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09342__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08145__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06388__I _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09893__A2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12751__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10988_ _05217_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09645__A2 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07656__A1 u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12727_ _01224_ net128 u_cpu.rf_ram.memory\[79\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06459__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11452__A2 _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12658_ _01155_ net241 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07012__I _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11204__A2 _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11609_ _00131_ net381 u_cpu.rf_ram.memory\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10007__A3 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout316_I net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12589_ _01087_ net172 u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__A1 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11469__I _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10963__A1 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__B1 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12131__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08908__A1 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08384__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ _03859_ _03877_ _03885_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06234__I2 u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06800__B _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12281__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05963_ _01604_ _01609_ _01611_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ u_cpu.rf_ram.memory\[72\]\[6\] _03836_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06490__S1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11849__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09333__A1 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07702_ _03154_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05894_ _01505_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08682_ u_cpu.rf_ram.memory\[141\]\[2\] _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11140__A1 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09884__A2 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07633_ u_cpu.rf_ram.memory\[42\]\[1\] _03107_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07895__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ u_cpu.rf_ram.memory\[7\]\[3\] _03060_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09636__A2 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09303_ _04192_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06515_ u_cpu.rf_ram.memory\[120\]\[4\] u_cpu.rf_ram.memory\[121\]\[4\] u_cpu.rf_ram.memory\[122\]\[4\]
+ u_cpu.rf_ram.memory\[123\]\[4\] _01606_ _01837_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07647__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07495_ _02959_ _03011_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06446_ u_cpu.rf_ram.memory\[72\]\[3\] u_cpu.rf_ram.memory\[73\]\[3\] u_cpu.rf_ram.memory\[74\]\[3\]
+ u_cpu.rf_ram.memory\[75\]\[3\] _01867_ _01732_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09234_ _04097_ _04141_ _04148_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08018__I _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09165_ _04088_ _04104_ _04107_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06377_ _01796_ _02022_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10484__S _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06870__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08116_ u_cpu.rf_ram.memory\[76\]\[2\] _03433_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08072__A1 u_cpu.rf_ram.memory\[77\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09096_ u_cpu.rf_ram.memory\[130\]\[5\] _04055_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10954__A1 u_cpu.rf_ram.memory\[104\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ u_cpu.rf_ram.memory\[139\]\[2\] _03388_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06622__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12624__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08375__A2 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _04686_ _04687_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06481__S1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08949_ u_cpu.rf_ram.memory\[49\]\[6\] _03962_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09324__A1 u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08127__A2 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11960_ _00482_ net24 u_cpu.rf_ram.memory\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _05315_ _05363_ _05366_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11891_ _00413_ net182 u_cpu.rf_ram.memory\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ _05324_ _05313_ _05325_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12004__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07638__A1 u_cpu.rf_ram.memory\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11434__A2 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ u_cpu.rf_ram.memory\[94\]\[7\] _05270_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12512_ _01013_ net255 u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12154__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06700__I3 u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12443_ _00944_ net249 u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11198__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08063__A1 u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12374_ _00875_ net479 u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10945__A1 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10193__I _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _05625_ _05620_ _05627_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06613__A2 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09982__I _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ u_cpu.rf_ram.memory\[86\]\[0\] _05584_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10207_ _04689_ _04872_ _04873_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11187_ _05538_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08598__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11370__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10138_ _04170_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06472__S1 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09315__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10069_ _04658_ _04704_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11122__A1 _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07007__I _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__I3 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout266_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09618__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05983__S0 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout433_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11425__A2 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06067__B _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06300_ _01616_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10484__I0 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ _02713_ _02837_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06152__I1 u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06231_ _01752_ _01878_ _01485_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11189__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07677__I _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08054__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ u_cpu.rf_ram.memory\[60\]\[1\] u_cpu.rf_ram.memory\[61\]\[1\] u_cpu.rf_ram.memory\[62\]\[1\]
+ u_cpu.rf_ram.memory\[63\]\[1\] _01617_ _01619_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12647__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06093_ _01692_ _01718_ _01741_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07801__A1 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _02705_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09554__A1 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08357__A2 _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12797__CLK net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09852_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _04557_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout81_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10164__A2 _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11361__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05925__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _03440_ _03454_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06758__I3 u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09783_ _04511_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10052__B _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06995_ u_cpu.cpu.state.init_done _02618_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08734_ _03647_ _03821_ _03830_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05946_ _01532_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05877_ u_cpu.rf_ram.memory\[20\]\[0\] u_cpu.rf_ram.memory\[21\]\[0\] u_cpu.rf_ram.memory\[22\]\[0\]
+ u_cpu.rf_ram.memory\[23\]\[0\] _01524_ _01525_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08665_ _03743_ _03783_ _03789_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _03025_ _03089_ _03096_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08596_ _03743_ _03732_ _03744_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06540__B2 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07547_ u_cpu.rf_ram.memory\[1\]\[7\] _03038_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11416__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07478_ u_cpu.rf_ram.memory\[18\]\[1\] _03000_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08293__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ u_cpu.rf_ram.memory\[126\]\[7\] _04127_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06429_ _01616_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06694__I2 u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10227__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08045__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ u_cpu.rf_ram.memory\[22\]\[4\] _04091_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08596__A2 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _04009_ _04040_ _04048_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11110_ _05488_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12090_ _00604_ net71 u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11041_ _05443_ _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09545__A1 u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06359__A1 _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11352__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07020__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06749__I3 u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12992_ _00051_ net521 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11943_ _00465_ net69 u_cpu.rf_ram.memory\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08520__A2 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11874_ _00396_ net185 u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06382__I1 u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11407__A2 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ u_cpu.rf_ram.memory\[28\]\[0\] _05313_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10756_ _05270_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07626__A4 _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06685__I2 u_cpu.rf_ram.memory\[110\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10687_ _02943_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12426_ _00927_ net49 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08036__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__A2 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12357_ _00858_ net423 u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06598__A1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11308_ _05564_ _05608_ _05615_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12288_ _00789_ net380 u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09536__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11239_ _05555_ _05571_ _05574_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10146__A2 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout383_I net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05800_ u_cpu.cpu.decode.co_mem_word _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06780_ u_cpu.rf_ram.memory\[120\]\[7\] u_cpu.rf_ram.memory\[121\]\[7\] u_cpu.rf_ram.memory\[122\]\[7\]
+ u_cpu.rf_ram.memory\[123\]\[7\] _01606_ _01608_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06770__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07960__I _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__A2 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _03649_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06522__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07401_ _02943_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10098__I _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08381_ _03570_ _03597_ _03602_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07263_ _02763_ _02822_ _02823_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06214_ _01710_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09002_ _03738_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08027__A1 u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ _02729_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10909__A1 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06145_ _01567_ _01791_ _01792_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09775__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06076_ _01502_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07250__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09527__A1 _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout502 net503 net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09904_ _03275_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout513 net514 net513 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout524 net538 net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11334__A1 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10137__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout535 net536 net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ u_arbiter.i_wb_cpu_rdt\[15\] _04546_ _04547_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ u_arbiter.i_wb_cpu_rdt\[0\] _04495_ _04497_ _02649_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06978_ u_cpu.rf_ram_if.rdata0\[5\] _02602_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06761__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08717_ _03819_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05929_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09697_ _04446_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08502__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08648_ u_cpu.rf_ram.memory\[15\]\[5\] _03775_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12812__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08579_ _03013_ _03595_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _04810_ _05160_ _05166_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11590_ _00112_ net189 u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10736__I _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _05123_ _05118_ u_cpu.cpu.ctrl.o_ibus_adr\[10\]
+ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12962__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _05078_
+ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09766__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12211_ _00725_ net294 u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06124__S0 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__A1 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12142_ _00656_ net52 u_cpu.rf_ram.memory\[133\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10471__I _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12073_ _00587_ net63 u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11325__A1 _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06170__B _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11024_ u_cpu.rf_ram.memory\[105\]\[3\] _05436_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06052__I0 u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06752__A1 _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12975_ _00032_ net515 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ _00448_ net86 u_cpu.rf_ram.memory\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12492__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05938__S0 _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _00379_ net99 u_cpu.rf_ram.memory\[65\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10439__I0 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10808_ _05212_ _05295_ _05302_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11788_ _00310_ net166 u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10064__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10646__I _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10064__B2 _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06658__I2 u_cpu.rf_ram.memory\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10739_ _05196_ _05259_ _05261_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout229_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08009__A1 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12409_ _00910_ net486 u_cpu.rf_ram.memory\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10367__A2 _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11564__A1 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09509__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07950_ _03222_ _03314_ _03321_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06080__B _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05794__A2 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06901_ _01444_ _02463_ _02539_ _01460_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07881_ net2 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09620_ _03256_ _03197_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07904__B _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06832_ u_cpu.cpu.bufreg2.i_cnt_done _02469_ _02470_ _02472_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_42_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07690__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09551_ _04342_ _04353_ _04359_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06763_ _02039_ _02404_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ u_cpu.rf_ram.memory\[56\]\[1\] _03683_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09482_ u_cpu.rf_ram.memory\[35\]\[3\] _04313_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06694_ u_cpu.rf_ram.memory\[112\]\[6\] u_cpu.rf_ram.memory\[113\]\[6\] u_cpu.rf_ram.memory\[114\]\[6\]
+ u_cpu.rf_ram.memory\[115\]\[6\] _02066_ _01631_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout44_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08433_ _02932_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12985__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08364_ _03575_ _03584_ _03591_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10055__A1 _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _02575_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08799__A2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08295_ _03505_ _03539_ _03546_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__S0 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _02763_ _02807_ _02809_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12215__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07177_ _02744_ _02738_ _02739_ _02751_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_121_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11555__A1 _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10358__A2 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06106__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01513_ _01775_ _01521_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12365__CLK net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06059_ u_cpu.rf_ram.memory\[80\]\[0\] u_cpu.rf_ram.memory\[81\]\[0\] u_cpu.rf_ram.memory\[82\]\[0\]
+ u_cpu.rf_ram.memory\[83\]\[0\] _01706_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout310 net311 net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout321 net333 net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout332 net333 net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout343 net347 net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_119_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout354 net369 net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout365 net366 net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout376 net377 net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08723__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout387 net392 net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09818_ _04538_ _04539_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout398 net407 net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08696__I _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06734__A1 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09749_ _04444_ _04472_ _04481_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12760_ _01257_ net208 u_cpu.rf_ram.memory\[83\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _00233_ net403 u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12691_ _01188_ net170 u_cpu.rf_ram.memory\[101\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06593__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11642_ _00164_ net163 u_cpu.rf_ram.memory\[78\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _03294_ _05783_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10524_ _02710_ _05108_ _05111_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09739__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12708__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10455_ _05069_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11546__A1 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10349__A2 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08411__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _04812_ _05023_ _05030_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__I0 u_cpu.rf_ram.memory\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12125_ _00639_ net258 u_cpu.rf_ram.memory\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12056_ _00570_ net9 u_cpu.rf_ram.memory\[71\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08714__A2 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _05411_ _05420_ _05427_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06725__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout179_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11882__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12958_ u_cpu.cpu.o_wen1 net280 u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10285__A1 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11909_ _00431_ net275 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12889_ _01386_ net507 u_cpu.rf_ram.memory\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__B2 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06584__S0 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12238__CLK net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout513_I net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10588__A2 _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ u_scanchain_local.module_data_in\[34\] u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _02686_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08080_ _03325_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07453__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12388__CLK net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11537__A1 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07205__A2 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A1 u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08953__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06803__I2 u_cpu.rf_ram.memory\[78\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08982_ _03932_ _03982_ _03987_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06964__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10760__A2 _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ u_cpu.rf_ram.memory\[16\]\[6\] _03306_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07864_ u_cpu.rf_ram.memory\[4\]\[0\] _03260_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__A1 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05933__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ u_cpu.rf_ram.memory\[8\]\[0\] _04390_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06815_ _02188_ _02456_ _01556_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07795_ _02914_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10060__B _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13013__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09534_ _04173_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06746_ u_cpu.rf_ram.memory\[12\]\[7\] u_cpu.rf_ram.memory\[13\]\[7\] u_cpu.rf_ram.memory\[14\]\[7\]
+ u_cpu.rf_ram.memory\[15\]\[7\] _01550_ _01553_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06319__I1 u_cpu.rf_ram.memory\[81\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10276__A1 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09130__A2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09465_ _04258_ _04297_ _04304_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07141__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06677_ _01926_ _02319_ _01929_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06575__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ _03623_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__A2 _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09396_ u_cpu.rf_ram.memory\[91\]\[3\] _04254_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09140__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08347_ _03579_ _03566_ _03580_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07444__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ _03509_ _03527_ _03535_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07229_ _02686_ _02794_ _02795_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07995__A3 _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11528__A1 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11755__CLK net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10240_ _04861_ _04901_ _04903_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10200__A1 _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10171_ _04842_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06955__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10751__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout151 net158 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout162 net231 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout173 net174 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout184 net185 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout195 net202 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10503__A2 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05843__I _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06183__A2 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12812_ _01309_ net125 u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12743_ _01240_ net143 u_cpu.rf_ram.memory\[106\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06566__S0 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12674_ _01171_ net50 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__A1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10019__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11625_ _00147_ net217 u_cpu.rf_ram.memory\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06891__B1 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12530__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A1 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07435__A2 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11556_ u_cpu.rf_ram.memory\[23\]\[5\] _05770_ _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10507_ _04812_ _05095_ _05102_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11487_ u_cpu.rf_ram.memory\[98\]\[1\] _05731_ _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11519__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10990__A2 _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _05047_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12680__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07199__A1 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10860__S _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ u_cpu.cpu.genblk3.csr.timer_irq_r _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12108_ _00622_ net282 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout296_I net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12039_ _00553_ net22 u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09360__A2 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__I3 u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout463_I net469 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07371__A1 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06600_ _02055_ _02243_ _02058_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ _03010_ _03070_ _03072_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12060__CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10258__A1 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06531_ _02169_ _02171_ _02173_ _02175_ _01858_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06557__S0 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ _02918_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _01992_ _02107_ _01556_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08871__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ u_cpu.rf_ram.memory\[67\]\[2\] _03486_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ _04115_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06393_ _01628_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ u_cpu.rf_ram.memory\[75\]\[0\] _03443_ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08623__A1 u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10834__I _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08063_ u_cpu.rf_ram.memory\[77\]\[0\] _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05928__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ _02612_ _02635_ _02633_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09179__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08926__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__A2 _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06401__A3 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08965_ u_cpu.rf_ram.memory\[136\]\[4\] _03974_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07916_ _03295_ _03300_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08896_ u_cpu.rf_ram.memory\[39\]\[2\] _03933_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12403__CLK net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ u_cpu.rf_ram.memory\[50\]\[2\] _03249_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06004__I3 u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07362__A1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08974__I _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ _03139_ _03199_ _03204_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09103__A2 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _04332_ _04334_ _04336_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06729_ _02362_ _02371_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12553__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06548__S0 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09448_ _04293_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08862__A1 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ _03272_ _02573_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11410_ u_cpu.rf_ram.memory\[26\]\[2\] _05686_ _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12390_ _00891_ net475 u_cpu.rf_ram.memory\[115\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11341_ _04228_ _02515_ _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05838__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06720__S0 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11272_ _05568_ _05584_ _05593_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13011_ _00072_ net531 u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10223_ _04689_ _04873_ _04886_ _04887_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08917__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06928__A1 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10154_ _04782_ _04825_ _04826_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09590__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07274__B _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10085_ _03278_ _04612_ _04766_ _04768_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_48_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12083__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10987_ _05413_ _05402_ _05414_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12726_ _01223_ net128 u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08853__A1 u_cpu.rf_ram.memory\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11920__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12657_ _01154_ net194 u_cpu.rf_ram.memory\[96\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ _00130_ net381 u_cpu.rf_ram.memory\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12588_ _01086_ net172 u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09802__B1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout211_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10412__A1 _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11539_ _03643_ _05755_ _05763_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout309_I net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08081__A2 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__S0 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12426__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06234__I3 u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _03749_ _03833_ _03840_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05962_ _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07701_ _03130_ _03153_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08681_ _03794_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07344__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _01541_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12576__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06778__S0 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11140__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07632_ _03010_ _03106_ _03108_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07895__A2 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07563_ _02921_ _03056_ _03061_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09097__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ _04158_ _04193_ _04196_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06514_ _01582_ _02158_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08844__A1 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07647__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07494_ _01591_ _02887_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09233_ u_cpu.rf_ram.memory\[125\]\[5\] _04144_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06445_ _01862_ _02090_ _01865_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ u_cpu.rf_ram.memory\[128\]\[1\] _04105_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06376_ u_cpu.rf_ram.memory\[36\]\[3\] u_cpu.rf_ram.memory\[37\]\[3\] u_cpu.rf_ram.memory\[38\]\[3\]
+ u_cpu.rf_ram.memory\[39\]\[3\] _01797_ _01586_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06458__I0 u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08115_ _03428_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10564__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__A2 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09095_ _04005_ _04051_ _04058_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06702__S0 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08046_ _03383_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05830__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09997_ _04655_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06386__A2 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _03939_ _03959_ _03966_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09324__A2 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08879_ u_cpu.rf_ram.memory\[138\]\[5\] _03918_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07335__A1 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06769__S0 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10910_ u_cpu.rf_ram.memory\[102\]\[1\] _05364_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11890_ _00412_ net270 u_cpu.rf_ram.memory\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11943__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05897__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10841_ u_cpu.rf_ram.memory\[28\]\[5\] _05318_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09088__A1 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _05218_ _05272_ _05280_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07638__A2 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08835__A1 _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12511_ _01012_ net183 u_cpu.rf_ram.memory\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06310__A2 _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12442_ _00943_ net249 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11198__A2 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A2 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12373_ _00874_ net479 u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07269__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__A2 _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06074__A1 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ u_cpu.rf_ram.memory\[88\]\[2\] _05626_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07810__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ _05582_ _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10206_ _04748_ _04782_ _04826_ _04793_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_49_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__A2 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11186_ _05538_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__A2 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12599__CLK net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06620__C _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10137_ _04812_ _04802_ _04813_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ _04726_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07326__A1 _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11122__A2 _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07877__A2 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout161_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout259_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__B _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05983__S1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07023__I _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12709_ _01206_ net135 u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout426_I net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07958__I _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06230_ u_cpu.rf_ram.memory\[132\]\[1\] u_cpu.rf_ram.memory\[133\]\[1\] u_cpu.rf_ram.memory\[134\]\[1\]
+ u_cpu.rf_ram.memory\[135\]\[1\] _01753_ _01754_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11189__A2 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06161_ _01799_ _01802_ _01804_ _01808_ _01613_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08054__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10936__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06092_ _01723_ _01729_ _01734_ _01739_ _01740_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07262__B1 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07801__A2 _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ _04609_ _04611_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11816__CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07693__I _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06811__B _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09851_ _04562_ _04563_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09554__A2 _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07565__A1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06612__I0 u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11361__A2 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08802_ _03861_ _03865_ _03874_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _04494_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06994_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] _02498_ u_cpu.cpu.state.o_cnt_r\[2\]
+ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11966__CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08733_ u_cpu.rf_ram.memory\[13\]\[7\] _03819_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05945_ u_cpu.rf_ram.memory\[32\]\[0\] u_cpu.rf_ram.memory\[33\]\[0\] u_cpu.rf_ram.memory\[34\]\[0\]
+ u_cpu.rf_ram.memory\[35\]\[0\] _01590_ _01593_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11113__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08664_ u_cpu.rf_ram.memory\[142\]\[3\] _03787_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05876_ _01506_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05941__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07615_ u_cpu.rf_ram.memory\[78\]\[4\] _03093_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ u_cpu.rf_ram.memory\[52\]\[3\] _03740_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__I2 u_cpu.rf_ram.memory\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _02946_ _03040_ _03048_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07477_ _02954_ _02999_ _03001_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08293__A2 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06143__I2 u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _04099_ _04129_ _04137_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06428_ _01494_ _02060_ _02073_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10227__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ _03745_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06359_ _01890_ _02004_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09078_ u_cpu.rf_ram.memory\[131\]\[6\] _04043_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ u_cpu.rf_ram.memory\[129\]\[3\] _03376_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11040_ _05404_ _05444_ _05447_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06359__A2 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11352__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10560__B1 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06012__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12991_ _00050_ net519 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11942_ _00464_ net71 u_cpu.rf_ram.memory\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05851__I _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ _00395_ net185 u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12121__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__A2 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06382__I2 u_cpu.rf_ram.memory\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10824_ _05311_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10615__A1 u_cpu.rf_ram.memory\[109\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10755_ _04295_ _03083_ _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09481__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10686_ _05215_ _05199_ _05216_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12425_ _00926_ net233 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08036__A2 _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11040__A1 _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12356_ _00857_ net472 u_cpu.rf_ram.memory\[121\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11307_ u_cpu.rf_ram.memory\[87\]\[5\] _05611_ _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12287_ _00788_ net400 u_cpu.rf_ram.memory\[91\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06631__B _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11989__CLK net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11238_ u_cpu.rf_ram.memory\[110\]\[1\] _05572_ _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09536__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11169_ u_cpu.rf_ram.memory\[59\]\[1\] _05527_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout376_I net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06522__A2 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06373__I2 u_cpu.rf_ram.memory\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ _02881_ u_cpu.rf_ram_if.wdata0_r\[6\] _02942_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_50_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ u_cpu.rf_ram.memory\[60\]\[2\] _03601_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12614__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07331_ u_cpu.cpu.decode.op26 _01449_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02880_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09472__A1 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08275__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07262_ _02808_ u_scanchain_local.module_data_in\[62\] _02788_ u_arbiter.i_wb_cpu_dbus_adr\[25\]
+ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__I3 u_cpu.rf_ram.memory\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09001_ _03998_ _03995_ _03999_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06213_ _01719_ _01860_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07193_ _02629_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08027__A2 _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12764__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11031__A1 _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06144_ _01520_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07786__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06075_ _01710_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05936__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _04444_ _04586_ _04595_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09527__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout503 net504 net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout514 net515 net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07538__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout525 net527 net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11334__A2 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout536 net537 net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _04544_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09765_ _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06977_ _01496_ _02591_ _02604_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__A2 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _03819_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11098__A1 u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05928_ _01576_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09696_ _04431_ _04447_ _04450_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08647_ _03638_ _03771_ _03778_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10845__A1 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10289__I _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ u_cpu.rf_ram.memory\[28\]\[0\] u_cpu.rf_ram.memory\[29\]\[0\] u_cpu.rf_ram.memory\[30\]\[0\]
+ u_cpu.rf_ram.memory\[31\]\[0\] _01504_ _01507_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A1 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12294__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08578_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ _02985_ _03037_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08266__A2 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07598__I _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__B _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__A1 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _05106_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10073__A2 _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ _02530_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12210_ _00724_ net300 u_cpu.rf_ram.memory\[126\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06007__I _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09766__A2 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11995__D _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06124__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12141_ _00655_ net43 u_cpu.rf_ram.memory\[133\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05846__I _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08222__I _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12072_ _00586_ net59 u_cpu.rf_ram.memory\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__A1 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11023_ _05406_ _05432_ _05437_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06201__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06052__I1 u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06752__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12974_ _00031_ net518 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12637__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10836__A1 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11925_ _00447_ net86 u_cpu.rf_ram.memory\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05938__S1 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11856_ _00378_ net98 u_cpu.rf_ram.memory\[65\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10807_ u_cpu.rf_ram.memory\[96\]\[4\] _05299_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10439__I1 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10927__I _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11661__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11787_ _00309_ net166 u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08257__A2 _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ u_cpu.rf_ram.memory\[97\]\[0\] _05260_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08009__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _05202_ _05198_ _05203_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12017__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12408_ _00909_ net486 u_cpu.rf_ram.memory\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11013__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10662__I _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12339_ _00840_ net477 u_cpu.rf_ram.memory\[120\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout493_I net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06900_ u_cpu.cpu.decode.co_ebreak _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _02952_ _03260_ _03269_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10524__B1 _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07971__I _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06831_ u_cpu.cpu.bufreg2.i_cnt_done u_cpu.cpu.immdec.imm31 _02471_ _02472_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06743__A2 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ u_cpu.rf_ram.memory\[120\]\[3\] _04357_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06762_ u_cpu.rf_ram.memory\[52\]\[7\] u_cpu.rf_ram.memory\[53\]\[7\] u_cpu.rf_ram.memory\[54\]\[7\]
+ u_cpu.rf_ram.memory\[55\]\[7\] _01647_ _02040_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08501_ _03661_ _03682_ _03684_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09481_ _04253_ _04309_ _04314_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06693_ _01660_ _02335_ _01611_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08496__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _03635_ _03624_ _03636_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout37_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10837__I _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ u_cpu.rf_ram.memory\[61\]\[4\] _03588_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09445__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _02513_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11252__A1 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10055__A2 _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ u_cpu.rf_ram.memory\[29\]\[4\] _03543_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06649__I3 u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07245_ _02808_ u_scanchain_local.module_data_in\[59\] _02788_ u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11004__A1 u_cpu.rf_ram.memory\[79\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07059__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _02751_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07759__A1 u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06106__S1 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11555__A2 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06127_ u_cpu.rf_ram.memory\[24\]\[1\] u_cpu.rf_ram.memory\[25\]\[1\] u_cpu.rf_ram.memory\[26\]\[1\]
+ u_cpu.rf_ram.memory\[27\]\[1\] _01516_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06431__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06058_ _01585_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout300 net302 net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout311 net312 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06982__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout322 net326 net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout333 net370 net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout344 net347 net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07881__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout355 net357 net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout366 net367 net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout377 net386 net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09817_ u_arbiter.i_wb_cpu_rdt\[10\] _04533_ _04534_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout388 net392 net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout399 net400 net399 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07931__A1 u_cpu.rf_ram.memory\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06734__A2 _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09748_ u_cpu.rf_ram.memory\[33\]\[7\] _04470_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__A1 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09679_ u_cpu.rf_ram.memory\[122\]\[4\] _04434_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11684__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__A2 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11710_ _00232_ net463 u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11491__A1 _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10294__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12690_ _01187_ net170 u_cpu.rf_ram.memory\[101\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09601__I _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06593__S1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11641_ _00163_ net163 u_cpu.rf_ram.memory\[78\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08239__A2 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09436__A1 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11243__A1 u_cpu.rf_ram.memory\[110\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11572_ _03279_ _05782_ _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07121__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10523_ _05113_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10597__A3 _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09739__A2 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _05066_
+ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11546__A2 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10385_ u_cpu.rf_ram.memory\[32\]\[4\] _05027_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08411__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _00638_ net258 u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12055_ _00569_ net9 u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07791__I _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11006_ u_cpu.rf_ram.memory\[79\]\[4\] _05424_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07922__A1 u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__S _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12957_ u_cpu.cpu.o_wen0 net279 u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06328__I2 u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11482__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11908_ _00430_ net275 u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12888_ _01385_ net506 u_cpu.rf_ram.memory\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06584__S1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout241_I net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09427__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11839_ _00361_ net97 u_cpu.rf_ram.memory\[67\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06356__B _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout339_I net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08650__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07966__I _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ u_arbiter.i_wb_cpu_rdt\[3\] _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__A3 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06413__A1 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08981_ u_cpu.rf_ram.memory\[135\]\[2\] _03986_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12802__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06964__A2 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07932_ _03224_ _03303_ _03310_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07407__S _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07863_ _03258_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__A2 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07913__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ _04388_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06814_ u_cpu.rf_ram.memory\[136\]\[7\] u_cpu.rf_ram.memory\[137\]\[7\] u_cpu.rf_ram.memory\[138\]\[7\]
+ u_cpu.rf_ram.memory\[139\]\[7\] _01759_ _02106_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12952__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07794_ _03210_ _03212_ _03214_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06110__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09533_ _04346_ _04335_ _04347_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06745_ _01547_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11473__A1 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ u_cpu.rf_ram.memory\[92\]\[4\] _04301_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06676_ u_cpu.rf_ram.memory\[48\]\[6\] u_cpu.rf_ram.memory\[49\]\[6\] u_cpu.rf_ram.memory\[50\]\[6\]
+ u_cpu.rf_ram.memory\[51\]\[6\] _01699_ _01927_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08415_ _03622_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06575__S1 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10567__I _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09395_ _04164_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_75_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08346_ u_cpu.rf_ram.memory\[62\]\[6\] _03571_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08277_ u_cpu.rf_ram.memory\[64\]\[6\] _03530_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07228_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _02783_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _02714_ _02736_ _02737_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12482__CLK net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10200__A2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _04599_ _04841_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06955__A2 _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout130 net141 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08157__A1 u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout141 net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout152 net158 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout163 net169 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout174 net178 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout185 net192 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10251__B _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06707__A2 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07904__A1 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout196 net201 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12811_ _01308_ net108 u_cpu.rf_ram.memory\[85\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06020__I _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10267__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12742_ _01239_ net143 u_cpu.rf_ram.memory\[106\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06566__S1 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A1 _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12673_ _01170_ net50 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08880__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11624_ _00146_ net217 u_cpu.rf_ram.memory\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10019__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _03637_ _05766_ _05773_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08632__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10506_ u_cpu.rf_ram.memory\[30\]\[4\] _05099_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11486_ _03620_ _05730_ _05732_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _05059_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08396__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _05018_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12107_ _00621_ net281 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10299_ u_cpu.cpu.immdec.imm19_12_20\[3\] _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08148__A1 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12038_ _00552_ net22 u_cpu.rf_ram.memory\[72\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout191_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08699__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout289_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__S0 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12205__CLK net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06530_ _02082_ _02174_ _02085_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11455__A1 _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06865__I u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10258__A2 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06557__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06461_ u_cpu.rf_ram.memory\[140\]\[3\] u_cpu.rf_ram.memory\[141\]\[3\] u_cpu.rf_ram.memory\[142\]\[3\]
+ u_cpu.rf_ram.memory\[143\]\[3\] _01993_ _02106_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06182__I0 u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08200_ _03481_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09180_ _04115_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06392_ _01622_ _02037_ _01626_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03441_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08623__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07696__I _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__B2 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ _03396_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10336__B _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ _02611_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08387__A1 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06105__I _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06937__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06788__I2 u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10850__I _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06493__S0 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08964_ _03935_ _03970_ _03976_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05944__I _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07915_ _01754_ _03297_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08895_ _03926_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__S0 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07846_ _03244_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07362__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07777_ u_cpu.rf_ram.memory\[43\]\[2\] _03203_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11446__A1 _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06728_ _02364_ _02366_ _02368_ _02370_ _01470_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09516_ u_cpu.rf_ram.memory\[117\]\[0\] _04335_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06548__S1 _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06708__C _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09447_ _04236_ u_cpu.cpu.state.o_cnt\[2\] _04233_ _00780_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06659_ _01468_ _02301_ _01521_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08862__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04244_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12848__CLK net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08329_ _03333_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09811__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11340_ _05636_ _05621_ _05637_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__S1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11271_ u_cpu.rf_ram.memory\[86\]\[7\] _05582_ _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12998__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10709__B1 _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13010_ _00071_ net530 u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08378__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10222_ _04722_ _04693_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06228__I1 u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10185__A1 _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06928__A2 _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _04634_ _04743_ _04764_ _04745_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_79_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05854__I _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07047__S _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _04617_ _04767_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__B2 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08550__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11437__A1 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05803__B u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10986_ u_cpu.rf_ram.memory\[99\]\[5\] _05407_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12725_ _01222_ net124 u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08853__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10000__I _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12656_ _01153_ net154 u_cpu.rf_ram.memory\[96\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11607_ _00129_ net379 u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12587_ _01085_ net319 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09802__B2 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11538_ u_cpu.rf_ram.memory\[89\]\[6\] _05758_ _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__B _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06711__S1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13003__CLK net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout204_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ _05717_ _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10871__S _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09030__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10176__A1 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10670__I _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07592__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05961_ _01483_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ _03152_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08680_ _03736_ _03795_ _03798_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05892_ _01540_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08541__A1 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07344__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07631_ u_cpu.rf_ram.memory\[42\]\[0\] _03107_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06778__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07562_ u_cpu.rf_ram.memory\[7\]\[2\] _03060_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11428__A1 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09097__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ u_cpu.rf_ram.memory\[38\]\[1\] _04194_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06513_ u_cpu.rf_ram.memory\[124\]\[4\] u_cpu.rf_ram.memory\[125\]\[4\] u_cpu.rf_ram.memory\[126\]\[4\]
+ u_cpu.rf_ram.memory\[127\]\[4\] _01947_ _01669_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07493_ _02907_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10100__A1 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08844__A2 _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _04095_ _04140_ _04147_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06444_ u_cpu.rf_ram.memory\[68\]\[3\] u_cpu.rf_ram.memory\[69\]\[3\] u_cpu.rf_ram.memory\[70\]\[3\]
+ u_cpu.rf_ram.memory\[71\]\[3\] _01725_ _01863_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10651__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09163_ _04083_ _04104_ _04106_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06375_ _02013_ _02015_ _02018_ _02020_ _01578_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11895__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08114_ _03413_ _03429_ _03432_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10403__A2 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09094_ u_cpu.rf_ram.memory\[130\]\[4\] _04055_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06702__S1 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07280__A1 _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08045_ _03334_ _03384_ _03387_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05830__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__A1 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__S0 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09996_ _04622_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08947_ u_cpu.rf_ram.memory\[49\]\[5\] _03962_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12520__CLK net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08878_ _03855_ _03914_ _03921_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__A1 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07335__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06769__S1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07829_ u_cpu.rf_ram.memory\[47\]\[3\] _03237_ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06719__B _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11419__A1 _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _05214_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05897__A2 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09088__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10771_ u_cpu.rf_ram.memory\[94\]\[6\] _05275_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12510_ _01011_ net188 u_cpu.rf_ram.memory\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10642__A2 _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11998__D _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06310__A3 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12441_ _00942_ net247 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13026__CLK net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12372_ _00873_ net417 u_cpu.rf_ram.memory\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11323_ _05619_ _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06074__A2 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11254_ _05582_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05821__A2 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11618__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _04693_ _04871_ _04608_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11185_ _05537_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10136_ u_cpu.rf_ram.memory\[114\]\[4\] _04808_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10067_ _02491_ _04699_ _04752_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06385__I0 u_cpu.rf_ram.memory\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10330__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09079__A2 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout154_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10866__S _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _05400_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10633__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12708_ _01205_ net134 u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout321_I net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12639_ _01136_ net145 u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout419_I net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06160_ _01604_ _01806_ _01807_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10397__A1 _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07262__A1 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _01577_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06696__S0 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10149__A1 _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09850_ u_arbiter.i_wb_cpu_rdt\[19\] _04559_ _04560_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07565__A2 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08801_ u_cpu.rf_ram.memory\[71\]\[7\] _03863_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09781_ _04510_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06993_ _02616_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08732_ _03644_ _03821_ _03829_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05944_ _01592_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout67_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08514__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12693__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08663_ _03739_ _03783_ _03788_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05875_ _01503_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06376__I0 u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10321__A1 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _03023_ _03089_ _03095_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08594_ _03742_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07214__I _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07545_ u_cpu.rf_ram.memory\[1\]\[6\] _03043_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08817__A2 _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10624__A2 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07476_ u_cpu.rf_ram.memory\[18\]\[0\] _03000_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09490__A2 _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _02062_ _02064_ _02068_ _02071_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09215_ u_cpu.rf_ram.memory\[126\]\[6\] _04132_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _04093_ _04085_ _04094_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12073__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06358_ u_cpu.rf_ram.memory\[20\]\[3\] u_cpu.rf_ram.memory\[21\]\[3\] u_cpu.rf_ram.memory\[22\]\[3\]
+ u_cpu.rf_ram.memory\[23\]\[3\] _01891_ _02003_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10388__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07253__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _04007_ _04040_ _04047_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06289_ _01646_ _01935_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08028_ _03337_ _03372_ _03377_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05803__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08753__A1 u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11910__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _04281_ _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12990_ _00049_ net519 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11941_ _00463_ net71 u_cpu.rf_ram.memory\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10312__A1 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _00394_ net183 u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07124__I _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10823_ _05311_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__A1 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10754_ _05221_ _05260_ _05269_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12416__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09481__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07492__A1 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10685_ u_cpu.rf_ram.memory\[93\]\[5\] _05206_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12424_ _00925_ net233 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10379__A1 _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09233__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11040__A2 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12355_ _00856_ net471 u_cpu.rf_ram.memory\[121\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08992__A1 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ _05562_ _05607_ _05614_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12286_ _00787_ net399 u_cpu.rf_ram.memory\[91\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _05550_ _05571_ _05573_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07547__A2 _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__A1 _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11168_ _05468_ _05526_ _05528_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10119_ _04151_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11099_ _05484_ _05471_ _05485_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout271_I net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10303__A1 _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout369_I net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06602__S0 _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07034__I u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06522__A3 _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout536_I net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07330_ _02876_ _02877_ _02878_ _02467_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__06873__I u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12096__CLK net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__A2 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07261_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _02818_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10082__A3 _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12909__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09000_ u_cpu.rf_ram.memory\[134\]\[1\] _03996_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06212_ u_cpu.rf_ram.memory\[64\]\[1\] u_cpu.rf_ram.memory\[65\]\[1\] u_cpu.rf_ram.memory\[66\]\[1\]
+ u_cpu.rf_ram.memory\[67\]\[1\] _01720_ _01721_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10328__C _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07192_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02753_ _02765_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09224__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06143_ u_cpu.rf_ram.memory\[12\]\[1\] u_cpu.rf_ram.memory\[13\]\[1\] u_cpu.rf_ram.memory\[14\]\[1\]
+ u_cpu.rf_ram.memory\[15\]\[1\] _01570_ _01572_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11031__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07786__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08983__A1 u_cpu.rf_ram.memory\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06074_ _01719_ _01722_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11933__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10790__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09902_ u_cpu.rf_ram.memory\[113\]\[7\] _04584_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout504 net508 net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout515 net518 net515 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07538__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08735__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout526 net527 net526 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout537 net538 net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09833_ _04549_ _04550_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _04494_ _04485_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06976_ u_cpu.rf_ram_if.rdata0\[4\] _02602_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05952__I _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ _03818_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05927_ _01486_ _01487_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09695_ u_cpu.rf_ram.memory\[115\]\[1\] _04448_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08646_ u_cpu.rf_ram.memory\[15\]\[4\] _03775_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05858_ _01506_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07710__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05789_ _01437_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08577_ _02905_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07528_ _03036_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ _02969_ _02987_ _02990_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11270__A2 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _05077_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09215__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07226__A1 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ u_cpu.rf_ram.memory\[12\]\[7\] _04064_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11022__A2 _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__A2 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12140_ _00654_ net53 u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10781__A1 _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12071_ _00585_ net59 u_cpu.rf_ram.memory\[143\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07529__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07119__I _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08726__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11022_ u_cpu.rf_ram.memory\[105\]\[2\] _05436_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06023__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06201__A2 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05862__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10701__C _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07055__S _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11089__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12973_ _00030_ net516 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09151__A1 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11924_ _00446_ net73 u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A2 _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11855_ _00377_ net97 u_cpu.rf_ram.memory\[65\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11806__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07789__I _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _05209_ _05295_ _05301_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05811__B _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11786_ _00308_ net268 u_cpu.rf_ram.memory\[139\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07465__A1 u_cpu.rf_ram.memory\[81\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10737_ _05258_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11261__A2 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11956__CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10668_ u_cpu.rf_ram.memory\[93\]\[1\] _05199_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12407_ _00908_ net485 u_cpu.rf_ram.memory\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07217__A1 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout117_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _03131_ _05158_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06642__B _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A1 u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08413__I _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12338_ _00839_ net365 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10772__A1 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A2 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12269_ _00770_ net358 u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__I0 u_cpu.rf_ram.memory\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout486_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09390__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A2 _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06830_ _01443_ u_cpu.cpu.branch_op u_cpu.cpu.csr_d_sel _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06761_ _01651_ _02402_ _01520_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__A1 u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08500_ u_cpu.rf_ram.memory\[56\]\[0\] _03683_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09480_ u_cpu.rf_ram.memory\[35\]\[2\] _04313_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06692_ u_cpu.rf_ram.memory\[120\]\[6\] u_cpu.rf_ram.memory\[121\]\[6\] u_cpu.rf_ram.memory\[122\]\[6\]
+ u_cpu.rf_ram.memory\[123\]\[6\] _01606_ _01608_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09693__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ u_cpu.rf_ram.memory\[5\]\[3\] _03632_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__I0 u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12731__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08362_ _03573_ _03584_ _03590_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ _02863_ _02547_ _02865_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07456__A1 u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08293_ _03503_ _03539_ _03545_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07244_ _02628_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07208__A1 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _02724_ _02748_ _02750_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07059__I1 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05947__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ _01517_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08323__I _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__B _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06271__C _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A2 _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06057_ _01616_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout301 net302 net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout312 net321 net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout323 net326 net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout334 net338 net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout345 net347 net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout356 net357 net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08184__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _04531_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout367 net368 net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout378 net379 net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06814__S0 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout389 net392 net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12261__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _04442_ _04472_ _04480_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06959_ _02474_ u_cpu.rf_ram.rdata\[4\] _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08993__I _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _04167_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08629_ u_cpu.rf_ram.memory\[9\]\[6\] _03762_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07695__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__A2 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06727__B _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11640_ _00162_ net166 u_cpu.rf_ram.memory\[78\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11979__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07402__I _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10249__B _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11571_ _02885_ u_cpu.rf_ram_if.rcnt\[1\] _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10522_ _02699_ _05108_ _05111_ _02710_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10453_ _05068_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05857__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06462__B _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08947__A1 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10384_ _04810_ _05023_ _05029_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10754__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06422__A2 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12123_ _00637_ net258 u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12054_ _00568_ net8 u_cpu.rf_ram.memory\[71\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08175__A2 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ _05409_ _05420_ _05426_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09064__I _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07922__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06281__S1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09124__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09999__I _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10809__A2 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12956_ u_cpu.cpu.o_wdata1 net334 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07135__B1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07686__A1 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11907_ _00429_ net375 u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11482__A2 _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12887_ _01384_ net499 u_cpu.rf_ram.memory\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11838_ _00360_ net97 u_cpu.rf_ram.memory\[67\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09427__A2 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07438__A1 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout234_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11769_ _00291_ net394 u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10993__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout401_I net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12134__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A1 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09239__I _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06413__A2 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08980_ _03981_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07931_ u_cpu.rf_ram.memory\[16\]\[5\] _03306_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07862_ _03258_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11170__A1 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ _04388_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07913__A2 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06813_ _01560_ _02454_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ u_cpu.rf_ram.memory\[48\]\[0\] _03213_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09115__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09532_ u_cpu.rf_ram.memory\[117\]\[5\] _04340_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06744_ u_cpu.rf_ram.memory\[8\]\[7\] u_cpu.rf_ram.memory\[9\]\[7\] u_cpu.rf_ram.memory\[10\]\[7\]
+ u_cpu.rf_ram.memory\[11\]\[7\] _02016_ _01507_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__I3 u_cpu.rf_ram.memory\[83\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ _04256_ _04297_ _04303_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06675_ _02039_ _02317_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11473__A2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__I0 u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06547__B _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08414_ _02961_ _03036_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09394_ _04253_ _04248_ _04255_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11225__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ _03349_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _03507_ _03527_ _03534_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10984__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07227_ _02703_ _02792_ _02793_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A1 u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _02721_ u_scanchain_local.module_data_in\[44\] _02722_ u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__12627__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ _01538_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07601__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07089_ u_arbiter.i_wb_cpu_rdt\[28\] u_arbiter.i_wb_cpu_dbus_dat\[25\] _02677_ _02682_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout120 net122 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout142 net162 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout153 net157 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12777__CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout164 net165 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06168__A1 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout175 net176 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11161__A1 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout186 net191 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10251__C _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout197 net201 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12810_ _01307_ net119 u_cpu.rf_ram.memory\[85\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12007__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09657__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12741_ _01238_ net115 u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06457__B _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12672_ _01169_ net49 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09409__A2 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07132__I _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A1 _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11623_ _00145_ net198 u_cpu.rf_ram.memory\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11216__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11554_ u_cpu.rf_ram.memory\[23\]\[4\] _05770_ _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10505_ _04810_ _05095_ _05101_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11485_ u_cpu.rf_ram.memory\[98\]\[0\] _05731_ _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10436_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _05054_
+ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08396__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09593__A1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08898__I _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10367_ u_cpu.cpu.immdec.imm31 _04670_ _04772_ _05016_ _05017_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_98_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12106_ _00620_ net273 u_cpu.rf_ram.memory\[137\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10298_ _04954_ _04948_ _04955_ _04752_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08148__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12037_ _00551_ net22 u_cpu.rf_ram.memory\[72\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__A2 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06254__S1 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout184_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10869__S _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07659__A1 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11455__A2 _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12939_ u_cpu.rf_ram_if.wdata0_r\[4\] net339 u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout351_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout449_I net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06706__I0 u_cpu.rf_ram.memory\[84\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08320__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06460_ _01721_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06391_ u_cpu.rf_ram.memory\[56\]\[3\] u_cpu.rf_ram.memory\[57\]\[3\] u_cpu.rf_ram.memory\[58\]\[3\]
+ u_cpu.rf_ram.memory\[59\]\[3\] _01623_ _01812_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08130_ _03441_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09820__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08061_ _03396_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06190__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07012_ _02633_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10718__A1 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11674__CLK net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08387__A2 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__A1 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout97_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__A1 _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08601__I _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ u_cpu.rf_ram.memory\[136\]\[3\] _03974_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06493__S1 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__A1 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08139__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07914_ _03299_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08894_ _03738_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09887__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06245__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07845_ _03215_ _03245_ _03248_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _03198_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09515_ _04333_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06727_ _01992_ _02369_ _01556_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11446__A2 _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08311__A2 _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09446_ _04280_ _04292_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06658_ u_cpu.rf_ram.memory\[12\]\[6\] u_cpu.rf_ram.memory\[13\]\[6\] u_cpu.rf_ram.memory\[14\]\[6\]
+ u_cpu.rf_ram.memory\[15\]\[6\] _01550_ _01553_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09377_ _04234_ u_cpu.cpu.state.o_cnt_r\[0\] _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_90_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06589_ _01926_ _02232_ _01929_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08075__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08328_ _03563_ _03565_ _03567_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10957__A1 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09811__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07822__A1 u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ u_cpu.rf_ram.memory\[65\]\[7\] _03513_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11270_ _05566_ _05584_ _05592_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10709__A1 _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10709__B2 _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09575__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08378__A2 _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _04672_ _04781_ _04871_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11382__A1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10185__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09607__I _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06928__A3 _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _04648_ _04726_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06484__S1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _04607_ _04732_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11134__A1 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__A2 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06031__I _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_2_539 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07063__S _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11437__A2 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10985_ _05214_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12724_ _01221_ net124 u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06313__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12655_ _01152_ net156 u_cpu.rf_ram.memory\[96\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11606_ _00128_ net379 u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08066__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12586_ _01084_ net319 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11697__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11537_ _03640_ _05755_ _05762_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07813__A1 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10156__C _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11468_ _02969_ _05718_ _05721_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09566__A1 _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08369__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _05048_
+ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11399_ _05634_ _05671_ _05679_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06650__B _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11373__A1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08421__I _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout399_I net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13039__I u_scanchain_local.data_out vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05960_ u_cpu.rf_ram.memory\[44\]\[0\] u_cpu.rf_ram.memory\[45\]\[0\] u_cpu.rf_ram.memory\[46\]\[0\]
+ u_cpu.rf_ram.memory\[47\]\[0\] _01606_ _01608_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09869__A2 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05891_ _01514_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12322__CLK net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07630_ _03105_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__I _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07895__A4 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07561_ _03055_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11428__A2 _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09300_ _04152_ _04193_ _04195_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06512_ _02150_ _02152_ _02154_ _02156_ _01832_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_55_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _02982_ _03000_ _03009_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06304__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__I1 u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10100__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12472__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09231_ u_cpu.rf_ram.memory\[125\]\[4\] _04144_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06443_ _01971_ _02088_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06374_ _01567_ _02019_ _01792_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09162_ u_cpu.rf_ram.memory\[128\]\[0\] _04105_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout12_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10939__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ u_cpu.rf_ram.memory\[76\]\[1\] _03430_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06607__A2 _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07804__A1 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ _04003_ _04051_ _04057_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06458__I2 u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10066__C _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06116__I _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08044_ u_cpu.rf_ram.memory\[139\]\[1\] _03385_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09557__A1 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07407__I1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05955__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10167__A2 _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07032__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09995_ _04649_ _04684_ _04665_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_88_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09309__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _03937_ _03958_ _03965_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11116__A1 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06791__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ u_cpu.rf_ram.memory\[138\]\[4\] _03918_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08532__A2 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07828_ _03217_ _03233_ _03238_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11419__A2 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07759_ u_cpu.rf_ram.memory\[41\]\[4\] _03189_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10770_ _05215_ _05272_ _05279_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _04264_ _04268_ _04277_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06846__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12440_ _00941_ net246 u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08048__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07410__I _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09796__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08599__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12371_ _00872_ net414 u_cpu.rf_ram.memory\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11322_ _02919_ _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__A1 u_cpu.rf_ram.memory\[120\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11253_ _05512_ _03453_ _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05865__I u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09337__I _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ _04638_ _04705_ _04690_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_10_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11184_ _03256_ _03102_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12345__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _04167_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11107__A1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10066_ _04740_ _04733_ _04741_ _04751_ _04676_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__09720__A1 u_cpu.rf_ram.memory\[116\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12495__CLK net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08287__A1 u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _05400_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12707_ _01204_ net171 u_cpu.rf_ram.memory\[103\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10899_ u_cpu.rf_ram.memory\[101\]\[5\] _05355_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08039__A1 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12638_ _01135_ net146 u_cpu.rf_ram.memory\[94\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__C _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09787__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout314_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12569_ _01067_ net323 u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10397__A2 _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06090_ _01735_ _01737_ _01738_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09539__A1 _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11346__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__A2 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09247__I _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06448__S1 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _03859_ _03865_ _03873_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A2 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06612__I2 u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ u_arbiter.i_wb_cpu_rdt\[2\] _04492_ _04509_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08731_ u_cpu.rf_ram.memory\[13\]\[6\] _03824_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05943_ _01591_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08514__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08662_ u_cpu.rf_ram.memory\[142\]\[2\] _03787_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05874_ _01467_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10321__A2 _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ u_cpu.rf_ram.memory\[78\]\[3\] _03093_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08593_ _02925_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11862__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12988__CLK net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07544_ _02940_ _03040_ _03047_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08278__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10085__A1 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06828__A2 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _02998_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09214_ _04097_ _04129_ _04136_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12218__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06426_ _01488_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08326__I _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09778__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ u_cpu.rf_ram.memory\[22\]\[3\] _04091_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06357_ _01736_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06288_ u_cpu.rf_ram.memory\[100\]\[2\] u_cpu.rf_ram.memory\[101\]\[2\] u_cpu.rf_ram.memory\[102\]\[2\]
+ u_cpu.rf_ram.memory\[103\]\[2\] _01934_ _01648_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09076_ u_cpu.rf_ram.memory\[131\]\[5\] _04043_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06687__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12368__CLK net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08027_ u_cpu.rf_ram.memory\[129\]\[2\] _03376_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11337__A1 _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__A1 _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08753__A2 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08996__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09978_ _04599_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08929_ u_cpu.rf_ram.memory\[137\]\[6\] _03950_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08505__A2 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11940_ _00462_ net68 u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06516__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10312__A2 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11871_ _00393_ net168 u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ _05310_ _03153_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11371__B _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10753_ u_cpu.rf_ram.memory\[97\]\[7\] _05258_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06819__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10871__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07492__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10684_ _05214_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12423_ _00924_ net234 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06127__S0 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12354_ _00855_ net362 u_cpu.rf_ram.memory\[121\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11305_ u_cpu.rf_ram.memory\[87\]\[4\] _05611_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12285_ _00786_ net400 u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11328__A1 _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11735__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11236_ u_cpu.rf_ram.memory\[110\]\[0\] _05572_ _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09941__A1 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ u_cpu.rf_ram.memory\[59\]\[0\] _05527_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _02499_ _04677_ _04799_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11098_ u_cpu.rf_ram.memory\[83\]\[6\] _05476_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10049_ _04625_ _04735_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__I1 u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10303__A2 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__S _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout264_I net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06602__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10067__A1 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10676__I _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout431_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout529_I net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10862__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07260_ _02817_ _02821_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07483__A2 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06286__A3 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08680__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06211_ _01849_ _01851_ _01854_ _01857_ _01858_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07191_ _02758_ _02753_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12510__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06142_ _01560_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08432__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06073_ u_cpu.rf_ram.memory\[64\]\[0\] u_cpu.rf_ram.memory\[65\]\[0\] u_cpu.rf_ram.memory\[66\]\[0\]
+ u_cpu.rf_ram.memory\[67\]\[0\] _01720_ _01721_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08983__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11300__I _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06994__A1 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10790__A2 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _04442_ _04586_ _04594_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12660__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout505 net506 net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout516 net517 net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout527 net529 net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09832_ u_arbiter.i_wb_cpu_rdt\[14\] _04546_ _04547_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08735__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout538 net1 net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06597__I1 u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09763_ _04494_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06975_ _01496_ _02589_ _02603_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13016__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _03050_ _03132_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05926_ _01567_ _01573_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09694_ _04425_ _04447_ _04449_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08645_ _03635_ _03771_ _03777_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05857_ _01505_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12040__CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08576_ _03679_ _03719_ _03728_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05788_ u_cpu.cpu.csr_imm _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07527_ _02870_ _02962_ _03035_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__11608__CLK net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10853__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ u_cpu.rf_ram.memory\[81\]\[1\] _02988_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08671__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06409_ _01659_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12190__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _02933_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__A1 u_cpu.rf_ram.memory\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _02951_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _04009_ _04028_ _04036_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10781__A2 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12070_ _00584_ net59 u_cpu.rf_ram.memory\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06037__I0 u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08726__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _05431_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09923__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06588__I1 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12972_ _00029_ net517 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11923_ _00445_ net73 u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11854_ _00376_ net99 u_cpu.rf_ram.memory\[65\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10049__A1 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ u_cpu.rf_ram.memory\[96\]\[3\] _05299_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11785_ _00307_ net274 u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12533__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10736_ _05258_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07465__A2 _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10667_ _05201_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12406_ _00907_ net465 u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08414__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12683__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _05157_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10221__A1 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12337_ _00838_ net365 u_cpu.rf_ram.memory\[120\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10772__A2 _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06214__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12268_ _00769_ net356 u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09914__A1 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ u_cpu.rf_ram.memory\[85\]\[3\] _05558_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12199_ _00713_ net343 u_cpu.rf_ram.memory\[127\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10524__A2 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__I _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__A2 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout381_I net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout479_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ u_cpu.rf_ram.memory\[56\]\[7\] u_cpu.rf_ram.memory\[57\]\[7\] u_cpu.rf_ram.memory\[58\]\[7\]
+ u_cpu.rf_ram.memory\[59\]\[7\] _01652_ _01552_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06691_ _01582_ _02333_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06200__I0 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ _03634_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__I _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08361_ u_cpu.rf_ram.memory\[61\]\[3\] _03588_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06339__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07312_ _02461_ _02864_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10339__C _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08653__A1 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ u_cpu.rf_ram.memory\[29\]\[3\] _03543_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11900__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _02804_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08405__A1 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ _02749_ u_scanchain_local.module_data_in\[47\] _02730_ u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10212__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ _01500_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08956__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__A1 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10763__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout302 net303 net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09905__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08708__A2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout313 net314 net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout324 net326 net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout335 net338 net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout346 net347 net346 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _04536_ _04537_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout357 net368 net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06814__S1 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout368 net369 net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout379 net385 net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07392__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ u_cpu.rf_ram.memory\[33\]\[6\] _04475_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06958_ _02584_ _02591_ _02592_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10279__A1 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05909_ _01510_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _04436_ _04428_ _04437_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _02527_ _01451_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12556__CLK net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _03641_ _03759_ _03766_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07695__A2 _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08892__A1 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08559_ _03717_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11205__I _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _05781_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09841__B1 _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10521_ _05112_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10452_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _05066_
+ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10383_ u_cpu.rf_ram.memory\[32\]\[3\] _05027_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06958__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10754__A2 _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12122_ _00636_ net265 u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06034__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12053_ _00567_ net8 u_cpu.rf_ram.memory\[71\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10506__A2 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11004_ u_cpu.rf_ram.memory\[79\]\[3\] _05424_ _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09372__A2 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06430__I0 u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09124__A2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12955_ u_cpu.rf_ram_if.wdata1_r\[7\] net335 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07135__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11906_ _00428_ net271 u_cpu.rf_ram.memory\[60\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12886_ _01383_ net497 u_cpu.rf_ram.memory\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07686__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A1 u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11923__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10690__A1 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11837_ _00359_ net97 u_cpu.rf_ram.memory\[67\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07438__A2 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11768_ _00290_ net394 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09832__B1 _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10719_ _03084_ _05233_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout227_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11699_ _00221_ net390 u_cpu.rf_ram.memory\[43\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10993__A2 _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__I _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10745__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12429__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07930_ _03222_ _03302_ _03309_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06879__I _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__I _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ _03257_ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09600_ _03037_ _03328_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12579__CLK net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11170__A2 _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06812_ u_cpu.rf_ram.memory\[140\]\[7\] u_cpu.rf_ram.memory\[141\]\[7\] u_cpu.rf_ram.memory\[142\]\[7\]
+ u_cpu.rf_ram.memory\[143\]\[7\] _01542_ _01544_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07792_ _03211_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09531_ _04170_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06743_ _01528_ _02384_ _01534_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ u_cpu.rf_ram.memory\[92\]\[3\] _04301_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout42_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08874__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06674_ u_cpu.rf_ram.memory\[52\]\[6\] u_cpu.rf_ram.memory\[53\]\[6\] u_cpu.rf_ram.memory\[54\]\[6\]
+ u_cpu.rf_ram.memory\[55\]\[6\] _01647_ _02040_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06724__I1 u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08413_ _03620_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ u_cpu.rf_ram.memory\[91\]\[2\] _04254_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08344_ _03577_ _03566_ _03578_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08626__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06119__I _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ u_cpu.rf_ram.memory\[64\]\[5\] _03530_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05958__I _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07226_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] u_cpu.cpu.ctrl.o_ibus_adr\[18\] _02765_ _02780_
+ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08929__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07157_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _02735_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09051__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06108_ _01752_ _01755_ _01756_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07088_ _02681_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07601__A2 _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06039_ _01683_ _01686_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout110 net123 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout132 net135 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09354__A2 _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout154 net157 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06168__A2 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout165 net169 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout176 net178 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11161__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__S0 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout187 net188 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10104__I _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout198 net200 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11946__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _04444_ _04460_ _04469_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06738__B _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12740_ _01237_ net115 u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A1 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07413__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06715__I1 u_cpu.rf_ram.memory\[77\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12671_ _01168_ net49 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A2 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11622_ _00144_ net209 u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06029__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06479__I0 u_cpu.rf_ram.memory\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11553_ _03634_ _05766_ _05772_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06473__B _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ u_cpu.rf_ram.memory\[30\]\[3\] _05099_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11484_ _05729_ _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10435_ _05058_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09042__A1 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10727__A2 _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09593__A2 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10366_ _04958_ _04911_ _04824_ _04717_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10723__B _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12105_ _00619_ net269 u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10297_ u_cpu.cpu.immdec.imm19_12_20\[3\] _04949_ _04952_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09345__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12036_ _00550_ net26 u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10014__I _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12871__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07108__A1 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout177_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08856__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07659__A2 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12938_ u_cpu.rf_ram_if.wdata0_r\[3\] net339 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12101__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12869_ _01366_ net496 u_cpu.rf_ram.memory\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06331__A2 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06182__I2 u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08608__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ _01919_ _02035_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09805__B1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10684__I _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout511_I net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08154__I _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ _03395_ _03132_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07831__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05842__A1 _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07011_ _02608_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06190__S1 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09033__A1 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10718__A2 _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__A2 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07595__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06398__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__A2 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08962_ _03932_ _03970_ _03975_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ _03279_ _03294_ _03297_ _03298_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11969__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09336__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08893_ _03930_ _03927_ _03931_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__A1 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07844_ u_cpu.rf_ram.memory\[50\]\[1\] _03246_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _03137_ _03199_ _03202_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06558__B _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09514_ _04333_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06726_ u_cpu.rf_ram.memory\[140\]\[6\] u_cpu.rf_ram.memory\[141\]\[6\] u_cpu.rf_ram.memory\[142\]\[6\]
+ u_cpu.rf_ram.memory\[143\]\[6\] _01993_ _02106_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08329__I _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10654__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _04281_ _04291_ _00773_ _02617_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06657_ _01547_ _02299_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A2 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09376_ _03271_ _02462_ _04240_ _04243_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06588_ u_cpu.rf_ram.memory\[48\]\[5\] u_cpu.rf_ram.memory\[49\]\[5\] u_cpu.rf_ram.memory\[50\]\[5\]
+ u_cpu.rf_ram.memory\[51\]\[5\] _01699_ _01927_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10406__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08327_ u_cpu.rf_ram.memory\[62\]\[0\] _03566_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08075__A2 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06293__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03509_ _03515_ _03523_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07822__A2 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__I _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08189_ _03424_ _03470_ _03478_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10709__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10220_ _04840_ _04885_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09575__A2 _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06228__I3 u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11382__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _04748_ _04823_ _04624_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_79_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10590__B1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__I _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12894__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ _04650_ _04763_ _04765_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07338__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11134__A2 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11374__B _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _05411_ _05401_ _05412_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07143__I _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10645__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12723_ _01220_ net153 u_cpu.rf_ram.memory\[99\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06313__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12654_ _01151_ net160 u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12274__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11605_ _00127_ net416 u_cpu.rf_ram.memory\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08066__A2 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12585_ _01083_ net319 u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11070__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11536_ u_cpu.rf_ram.memory\[89\]\[5\] _05758_ _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07813__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10009__I _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11467_ u_cpu.rf_ram.memory\[0\]\[1\] _05719_ _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10418_ _05049_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09566__A2 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11398_ u_cpu.rf_ram.memory\[27\]\[6\] _05674_ _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _04774_ u_arbiter.i_wb_cpu_rdt\[18\] _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07318__I _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout294_I net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12019_ _00533_ net57 u_cpu.rf_ram.memory\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05890_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout461_I net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10679__I _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07560_ _02915_ _03056_ _03059_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08829__A1 u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12617__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10636__A1 _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06511_ _02055_ _02155_ _02058_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07491_ u_cpu.rf_ram.memory\[18\]\[7\] _02998_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07501__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06304__A2 _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04093_ _04140_ _04146_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ u_cpu.rf_ram.memory\[64\]\[3\] u_cpu.rf_ram.memory\[65\]\[3\] u_cpu.rf_ram.memory\[66\]\[3\]
+ u_cpu.rf_ram.memory\[67\]\[3\] _01720_ _01972_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ _04103_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06373_ u_cpu.rf_ram.memory\[12\]\[3\] u_cpu.rf_ram.memory\[13\]\[3\] u_cpu.rf_ram.memory\[14\]\[3\]
+ u_cpu.rf_ram.memory\[15\]\[3\] _01570_ _01572_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11641__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09254__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10939__A2 _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10347__C _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ _03408_ _03429_ _03431_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11061__A1 _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07002__B _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09092_ u_cpu.rf_ram.memory\[130\]\[3\] _04055_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07804__A2 _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__I3 u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05815__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08043_ _03326_ _03384_ _03386_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11791__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09994_ _04653_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10572__B1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ u_cpu.rf_ram.memory\[49\]\[4\] _03962_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11116__A2 _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08876_ _03853_ _03914_ _03920_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07040__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ u_cpu.rf_ram.memory\[47\]\[2\] _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10875__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07740__A1 u_cpu.rf_ram.memory\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07758_ _03142_ _03185_ _03191_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08059__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12297__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06709_ u_cpu.rf_ram.memory\[64\]\[6\] u_cpu.rf_ram.memory\[65\]\[6\] u_cpu.rf_ram.memory\[66\]\[6\]
+ u_cpu.rf_ram.memory\[67\]\[6\] _01731_ _01972_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10478__I1 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _03144_ _03134_ _03145_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08296__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09428_ u_cpu.rf_ram.memory\[90\]\[7\] _04266_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ _04230_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09245__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11052__A1 u_cpu.rf_ram.memory\[106\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12370_ _00871_ net423 u_cpu.rf_ram.memory\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11321_ _05623_ _05620_ _05624_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11252_ _05568_ _05572_ _05581_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09548__A2 _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ _04869_ _04870_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11183_ _05486_ _05527_ _05536_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08220__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10134_ _04810_ _04802_ _04811_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11107__A2 _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10065_ _04746_ _04750_ _04701_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05881__I _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07074__S _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10720__C _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__A1 _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09484__A1 u_cpu.rf_ram.memory\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10967_ _03166_ _05374_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08287__A2 _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12706_ _01203_ net137 u_cpu.rf_ram.memory\[103\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10898_ _05322_ _05351_ _05358_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05896__I1 u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12637_ _01134_ net152 u_cpu.rf_ram.memory\[94\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09236__A1 _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08039__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07098__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11043__A1 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06217__I _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12568_ _01066_ net323 u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11519_ _03643_ _05743_ _05751_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12499_ _01000_ net493 u_cpu.rf_ram.memory\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout307_I net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09528__I _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11346__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__A2 _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _02518_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _03641_ _03821_ _03828_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05942_ u_cpu.raddr\[1\] _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__I _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _03782_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05873_ _01513_ _01519_ _01521_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07722__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _03020_ _03089_ _03094_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ _03739_ _03732_ _03741_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10609__A1 u_cpu.rf_ram.memory\[109\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ u_cpu.rf_ram.memory\[1\]\[5\] _03043_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08278__A2 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__A1 _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10085__A2 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07474_ _02998_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06828__A3 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ u_cpu.rf_ram.memory\[126\]\[5\] _04132_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ _01683_ _02070_ _01687_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10077__C _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11034__A1 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07089__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09144_ _03742_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06356_ _01513_ _02000_ _02001_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09075_ _04005_ _04039_ _04046_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ _01568_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05966__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08026_ _03371_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08342__I _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11337__A2 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06213__A1 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__A2 _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09977_ _04608_ _04620_ _04625_ _04643_ _04668_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07961__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08928_ _03939_ _03947_ _03954_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10848__A1 _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09702__A2 _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08859_ u_cpu.rf_ram.memory\[14\]\[5\] _03906_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11687__CLK net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11208__I _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06516__A2 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12932__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11870_ _00392_ net183 u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _02963_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09466__A1 u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08269__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ _05218_ _05260_ _05268_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11273__A1 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10683_ _02937_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09218__A1 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11025__A1 _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12422_ _00923_ net234 u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09769__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06127__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10782__I _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12353_ _00854_ net364 u_cpu.rf_ram.memory\[121\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05876__I _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11304_ _05560_ _05607_ _05613_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12284_ _00785_ net399 u_cpu.rf_ram.memory\[91\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11235_ _05570_ _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12462__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__A2 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _05525_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _04740_ _04789_ _04798_ _04698_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_96_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11097_ _05217_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10839__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10048_ _04702_ _04730_ _04734_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06507__A2 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11500__A2 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__I2 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__I _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__A1 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout257_I net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11999_ _00004_ net291 u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11264__A1 _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__B _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06375__C _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout424_I net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08680__A2 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _01488_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06691__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ _02704_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ u_cpu.rf_ram.memory\[8\]\[1\] u_cpu.rf_ram.memory\[9\]\[1\] u_cpu.rf_ram.memory\[10\]\[1\]
+ u_cpu.rf_ram.memory\[11\]\[1\] _01561_ _01564_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10692__I _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08432__A2 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05786__I _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05877__S0 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06072_ _01505_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12805__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06994__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09900_ u_cpu.rf_ram.memory\[113\]\[6\] _04589_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout506 net507 net506 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout517 net518 net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09831_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _04544_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09932__A2 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout528 net529 net528 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07943__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06597__I2 u_cpu.rf_ram.memory\[110\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09762_ _02632_ _02622_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06974_ u_cpu.rf_ram_if.rdata0\[3\] _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout72_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10360__C _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06410__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05925_ _01484_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08713_ _03755_ _03808_ _03817_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09693_ u_cpu.rf_ram.memory\[115\]\[0\] _04448_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09696__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08644_ u_cpu.rf_ram.memory\[15\]\[3\] _03775_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05856_ u_cpu.raddr\[1\] _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ u_cpu.rf_ram.memory\[53\]\[7\] _03717_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05787_ _01438_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ _03033_ _02892_ _03034_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__B _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07457_ _02954_ _02987_ _02989_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12335__CLK net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08671__A2 _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06682__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06408_ _01941_ _02053_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11007__A1 _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07388_ _02932_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11558__A2 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09127_ _04079_ _04066_ _04080_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06339_ u_cpu.rf_ram.memory\[136\]\[2\] u_cpu.rf_ram.memory\[137\]\[2\] u_cpu.rf_ram.memory\[138\]\[2\]
+ u_cpu.rf_ram.memory\[139\]\[2\] _01747_ _01875_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08423__A2 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09620__A1 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07226__A3 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12485__CLK net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ u_cpu.rf_ram.memory\[132\]\[6\] _04031_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08009_ u_cpu.rf_ram.memory\[119\]\[4\] _03362_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ _05404_ _05432_ _05435_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09923__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07934__A1 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12971_ _00028_ net517 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11494__A1 u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11922_ _00444_ net213 u_cpu.rf_ram.memory\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10297__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10777__I _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ _00375_ net97 u_cpu.rf_ram.memory\[65\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__I2 u_cpu.rf_ram.memory\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10804_ _05205_ _05295_ _05300_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11246__A1 _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11784_ _00306_ net274 u_cpu.rf_ram.memory\[139\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08111__A1 u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _02984_ _05158_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08662__A2 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06673__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10666_ _02912_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12828__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11702__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12405_ _00906_ net485 u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09611__A1 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08414__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ u_cpu.cpu.immdec.imm11_7\[2\] _02897_ _03085_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_51_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05859__S0 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12336_ _00837_ net365 u_cpu.rf_ram.memory\[120\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06976__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12267_ _00768_ net356 u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12978__CLK net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08178__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11218_ _05208_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12198_ _00712_ net298 u_cpu.rf_ram.memory\[127\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07925__A1 u_cpu.rf_ram.memory\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__I2 u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11149_ u_cpu.rf_ram.memory\[84\]\[1\] _05515_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06690_ u_cpu.rf_ram.memory\[124\]\[6\] u_cpu.rf_ram.memory\[125\]\[6\] u_cpu.rf_ram.memory\[126\]\[6\]
+ u_cpu.rf_ram.memory\[127\]\[6\] _01947_ _01707_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09541__I _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08350__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10687__I _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11237__A1 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ _03570_ _03584_ _03589_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07311_ _02519_ _02525_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06339__S1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08291_ _03500_ _03539_ _03544_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09850__A1 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07996__I _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A1 _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ _02803_ _02805_ _02806_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07173_ _02628_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06124_ u_cpu.rf_ram.memory\[28\]\[1\] u_cpu.rf_ram.memory\[29\]\[1\] u_cpu.rf_ram.memory\[30\]\[1\]
+ u_cpu.rf_ram.memory\[31\]\[1\] _01504_ _01771_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09917__S _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06967__A2 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ _01558_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A1 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08620__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__A2 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout303 net304 net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout314 net320 net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout325 net326 net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout336 net337 net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_119_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09814_ u_arbiter.i_wb_cpu_rdt\[9\] _04533_ _04534_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xfanout347 net353 net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06275__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout358 net363 net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout369 net370 net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07236__I u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09745_ _04440_ _04472_ _04479_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09669__A1 u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06957_ _02587_ u_cpu.rf_ram_if.rdata1\[3\] _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05908_ _01547_ _01554_ _01556_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ u_cpu.rf_ram.memory\[122\]\[3\] _04434_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06888_ _01443_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09451__I _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A1 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08627_ u_cpu.rf_ram.memory\[9\]\[5\] _03762_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05839_ _01489_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__I2 u_cpu.rf_ram.memory\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08558_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07509_ _02927_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08489_ u_cpu.rf_ram.memory\[57\]\[5\] _03669_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08644__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09841__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10520_ _02513_ _05108_ _05111_ _02699_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _05067_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11875__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11221__I _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10382_ _04807_ _05023_ _05028_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06958__A2 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12121_ _00635_ net274 u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12052_ _00566_ net9 u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11003_ _05406_ _05420_ _05425_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__S0 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07383__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06050__I _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12500__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12954_ u_cpu.rf_ram_if.wdata1_r\[6\] net335 u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11905_ _00427_ net271 u_cpu.rf_ram.memory\[60\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12885_ _01382_ net497 u_cpu.rf_ram.memory\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10690__A2 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11836_ _00358_ net105 u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12650__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09832__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11767_ _00289_ net345 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06646__A1 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _04674_ _05241_ _05243_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_35_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11698_ _00220_ net453 u_cpu.rf_ram.memory\[43\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout122_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ u_cpu.rf_ram.memory\[2\]\[3\] _05188_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09060__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__A2 u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12319_ _00820_ net488 u_cpu.rf_ram.memory\[34\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout491_I net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09899__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06257__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07860_ _03013_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06811_ _01763_ _02452_ _01485_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ _03211_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12180__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06742_ u_cpu.rf_ram.memory\[0\]\[7\] u_cpu.rf_ram.memory\[1\]\[7\] u_cpu.rf_ram.memory\[2\]\[7\]
+ u_cpu.rf_ram.memory\[3\]\[7\] _01529_ _01530_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09530_ _04344_ _04334_ _04345_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11748__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09271__I _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09461_ _04253_ _04297_ _04302_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06673_ _01651_ _02315_ _01520_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06724__I2 u_cpu.rf_ram.memory\[138\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ _02906_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10681__A2 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09392_ _04247_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08343_ u_cpu.rf_ram.memory\[62\]\[5\] _03571_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11898__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__B2 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06637__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06488__I1 u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _03505_ _03526_ _03533_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08615__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10366__B _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06563__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ _02790_ _02781_ _02791_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__I _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05860__A2 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _02725_ _02727_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09051__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06107_ _01533_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07087_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_dbus_dat\[24\] _02677_ _02681_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05974__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06038_ _01595_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout100 net103 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout111 net114 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout122 net123 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout133 net135 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__12523__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout144 net145 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout155 net156 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout166 net168 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout177 net178 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06799__S1 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout188 net191 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07989_ u_cpu.rf_ram.memory\[40\]\[6\] _03338_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ u_cpu.rf_ram.memory\[116\]\[7\] _04458_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08314__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09659_ u_cpu.rf_ram.memory\[112\]\[7\] _04413_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06715__I2 u_cpu.rf_ram.memory\[78\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06876__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12670_ _01167_ net48 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11621_ _00143_ net432 u_cpu.rf_ram.memory\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13029__CLK net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09814__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06628__A1 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06479__I1 u_cpu.rf_ram.memory\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11552_ u_cpu.rf_ram.memory\[23\]\[3\] _05770_ _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10503_ _04807_ _05095_ _05100_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11483_ _05729_ _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10434_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _05054_
+ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06045__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10188__A1 _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09042__A2 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10365_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _02715_ _05016_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05884__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09356__I _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06800__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12104_ _00618_ net273 u_cpu.rf_ram.memory\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ u_cpu.cpu.immdec.imm19_12_20\[2\] _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06239__S0 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12035_ _00549_ net24 u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08553__A1 u_cpu.rf_ram.memory\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__A2 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10360__A1 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10112__A1 _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12937_ u_cpu.rf_ram_if.wdata0_r\[2\] net340 u_cpu.rf_ram_if.wdata0_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08856__A2 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__A1 _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12868_ _01365_ net501 u_cpu.rf_ram.memory\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06182__I3 u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11819_ _00341_ net199 u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09805__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout337_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08608__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12799_ _01296_ net413 u_cpu.rf_ram.memory\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06664__B _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09805__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout504_I net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07010_ u_arbiter.i_wb_cpu_ack _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05842__A2 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09033__A2 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10179__B2 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07595__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08792__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08961_ u_cpu.rf_ram.memory\[136\]\[2\] _03974_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _01753_ _03296_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08892_ u_cpu.rf_ram.memory\[39\]\[1\] _03928_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _03210_ _03245_ _03247_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10351__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ u_cpu.rf_ram.memory\[43\]\[1\] _03200_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09513_ _02960_ _04179_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06725_ _01539_ _02367_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06158__I0 u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11036__I _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10654__A2 _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06656_ u_cpu.rf_ram.memory\[8\]\[6\] u_cpu.rf_ram.memory\[9\]\[6\] u_cpu.rf_ram.memory\[10\]\[6\]
+ u_cpu.rf_ram.memory\[11\]\[6\] _02016_ _01507_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06402__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09444_ _02493_ _04290_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09375_ _02498_ _04242_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06587_ _02039_ _02230_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05969__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12076__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10406__A2 _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08345__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _03564_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ u_cpu.rf_ram.memory\[65\]\[6\] _03518_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07208_ _02696_ _02776_ _02777_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08188_ u_cpu.rf_ram.memory\[68\]\[6\] _03473_ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07139_ _02608_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07586__A2 _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08783__A1 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _04822_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08080__I _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11913__CLK net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10081_ _04764_ _04643_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09904__I _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__A1 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10983_ u_cpu.rf_ram.memory\[99\]\[4\] _05407_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08838__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12722_ _01219_ net153 u_cpu.rf_ram.memory\[99\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06849__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10645__A2 _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12653_ _01150_ net205 u_cpu.rf_ram.memory\[96\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05879__I _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11604_ _00126_ net416 u_cpu.rf_ram.memory\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12584_ _01082_ net327 u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11070__A2 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11535_ _03637_ _05754_ _05761_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _02954_ _05718_ _05720_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07026__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10417_ u_arbiter.i_wb_cpu_dbus_adr\[2\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _05048_
+ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11397_ _05632_ _05671_ _05678_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11593__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10348_ _04753_ _04902_ _04998_ _05000_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10025__I _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _04938_ _04939_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07329__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__A1 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12018_ _00532_ net69 u_cpu.rf_ram.memory\[141\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10333__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout287_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06659__B _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06632__S0 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout454_I net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06510_ u_cpu.rf_ram.memory\[104\]\[4\] u_cpu.rf_ram.memory\[105\]\[4\] u_cpu.rf_ram.memory\[106\]\[4\]
+ u_cpu.rf_ram.memory\[107\]\[4\] _02056_ _01624_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12099__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10636__A2 _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07490_ _02980_ _03000_ _03008_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07501__A2 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06441_ _02077_ _02079_ _02081_ _02086_ _01858_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_61_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05789__I _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09160_ _04103_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06372_ _01560_ _02017_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ u_cpu.rf_ram.memory\[76\]\[0\] _03430_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09091_ _04000_ _04051_ _04056_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06312__I0 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11061__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ u_cpu.rf_ram.memory\[139\]\[0\] _03385_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05815__A2 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11936__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07509__I _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09993_ _04682_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06240__A2 _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08944_ _03935_ _03958_ _03964_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08517__A1 _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10324__A1 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08875_ u_cpu.rf_ram.memory\[138\]\[3\] _03918_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09190__A1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ _03232_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07040__I1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__S0 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ u_cpu.rf_ram.memory\[41\]\[3\] _03189_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10627__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06708_ _02344_ _02346_ _02348_ _02350_ _01689_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07688_ u_cpu.rf_ram.memory\[45\]\[4\] _03140_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04262_ _04268_ _04276_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06639_ _01992_ _02282_ _01574_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12711__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _03270_ _04229_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08309_ _03498_ _03552_ _03555_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11052__A2 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__I0 u_cpu.rf_ram.memory\[120\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09289_ _04168_ _04181_ _04188_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11320_ u_cpu.rf_ram.memory\[88\]\[1\] _05621_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__A1 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11251_ u_cpu.rf_ram.memory\[110\]\[7\] _05570_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08756__A1 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ u_cpu.cpu.immdec.imm24_20\[4\] _04842_ _04844_ u_cpu.cpu.immdec.imm30_25\[0\]
+ _04866_ _04772_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11182_ u_cpu.rf_ram.memory\[59\]\[7\] _05525_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ u_cpu.rf_ram.memory\[114\]\[3\] _04808_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08508__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10064_ _04748_ _04749_ _04642_ _04660_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06614__S0 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__I0 u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11809__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06993__I _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10966_ _05195_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09484__A2 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12705_ _01202_ net137 u_cpu.rf_ram.memory\[103\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06926__C _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12391__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11404__I _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10897_ u_cpu.rf_ram.memory\[101\]\[4\] _05355_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12636_ _01133_ net146 u_cpu.rf_ram.memory\[94\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09236__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__A2 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07098__I1 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12567_ _01065_ net310 u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__I _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11518_ u_cpu.rf_ram.memory\[100\]\[6\] _05746_ _05751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12498_ _00999_ net492 u_cpu.rf_ram.memory\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout202_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11449_ _05705_ _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08747__A1 u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11346__A3 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ _02524_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05941_ _01548_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05872_ _01520_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08660_ _03736_ _03783_ _03786_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07722__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07611_ u_cpu.rf_ram.memory\[78\]\[2\] _03093_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06376__I3 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08591_ u_cpu.rf_ram.memory\[52\]\[2\] _03740_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__B1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12734__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07542_ _02934_ _03039_ _03046_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09475__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _02891_ _02964_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09212_ _04095_ _04128_ _04135_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06424_ u_cpu.rf_ram.memory\[116\]\[3\] u_cpu.rf_ram.memory\[117\]\[3\] u_cpu.rf_ram.memory\[118\]\[3\]
+ u_cpu.rf_ram.memory\[119\]\[3\] _02069_ _01685_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09227__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11034__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06355_ _01484_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09143_ _04090_ _04085_ _04092_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07089__I1 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08986__A1 _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09074_ u_cpu.rf_ram.memory\[131\]\[4\] _04043_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06286_ _01499_ _01896_ _01908_ _01932_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ _03334_ _03372_ _03375_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08738__A1 u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06213__A2 _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ _04649_ _04667_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05982__I _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12264__CLK net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07961__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08927_ u_cpu.rf_ram.memory\[137\]\[5\] _03950_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05972__A1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09163__A1 _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _03638_ _03902_ _03909_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07174__B1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07713__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ u_cpu.rf_ram.memory\[48\]\[5\] _03218_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _03848_ _03864_ _03867_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10820_ _05195_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07477__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ u_cpu.rf_ram.memory\[97\]\[6\] _05263_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11273__A2 _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11224__I _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06318__I _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _05212_ _05198_ _05213_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09218__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _00922_ net235 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07229__A1 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11025__A2 _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08977__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12352_ _00853_ net364 u_cpu.rf_ram.memory\[121\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10784__A1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11303_ u_cpu.rf_ram.memory\[87\]\[3\] _05611_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12283_ _00784_ net398 u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__I _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12607__CLK net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11234_ _05570_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06053__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06988__I u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11165_ _05525_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05892__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07085__S _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _04791_ _04792_ _04797_ _04739_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11096_ _05482_ _05471_ _05483_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05963__A1 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09154__A1 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10047_ _04607_ _04642_ _04732_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07165__B1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__I3 u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11781__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11998_ _00003_ net295 u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout152_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ u_cpu.rf_ram.memory\[104\]\[0\] _05389_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11264__A2 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12619_ _01116_ net146 u_cpu.rf_ram.memory\[93\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout417_I net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ _01785_ _01787_ _01556_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08968__A1 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11567__A3 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10775__A1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01540_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06443__A2 _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05877__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12287__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06994__A3 _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08196__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout507 net508 net507 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09830_ _04545_ _04548_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout518 net524 net518 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout529 net537 net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_28_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ _02651_ _04490_ _04492_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06973_ _01471_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09145__A1 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ u_cpu.rf_ram.memory\[140\]\[7\] _03806_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05924_ u_cpu.rf_ram.memory\[12\]\[0\] u_cpu.rf_ram.memory\[13\]\[0\] u_cpu.rf_ram.memory\[14\]\[0\]
+ u_cpu.rf_ram.memory\[15\]\[0\] _01570_ _01572_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09692_ _04446_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09696__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08643_ _03631_ _03771_ _03776_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05855_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_81_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ _03677_ _03719_ _03727_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05786_ _01437_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07459__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ u_cpu.cpu.immdec.imm11_7\[3\] _02878_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06506__I0 u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06138__I _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ u_cpu.rf_ram.memory\[81\]\[0\] _02988_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06407_ u_cpu.rf_ram.memory\[108\]\[3\] u_cpu.rf_ram.memory\[109\]\[3\] u_cpu.rf_ram.memory\[110\]\[3\]
+ u_cpu.rf_ram.memory\[111\]\[3\] _02052_ _01827_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11007__A2 _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _02931_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05977__I _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08959__A1 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ u_cpu.rf_ram.memory\[12\]\[6\] _04071_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06338_ _01957_ _01984_ _01743_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__I _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10766__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09620__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06269_ u_cpu.rf_ram.memory\[44\]\[2\] u_cpu.rf_ram.memory\[45\]\[2\] u_cpu.rf_ram.memory\[46\]\[2\]
+ u_cpu.rf_ram.memory\[47\]\[2\] _01805_ _01608_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09057_ _04007_ _04028_ _04035_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _03341_ _03358_ _03364_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11654__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08187__A2 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05926__B _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06198__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07934__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__I3 u_cpu.rf_ram.memory\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ _04602_ _02642_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A1 _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12970_ _00027_ net517 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09912__I _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _00443_ net220 u_cpu.rf_ram.memory\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07698__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11494__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _00374_ net107 u_cpu.rf_ram.memory\[65\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07432__I _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ u_cpu.rf_ram.memory\[96\]\[2\] _05299_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11246__A2 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _00305_ net273 u_cpu.rf_ram.memory\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08111__A2 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ _02894_ _05224_ _05256_ _05257_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07870__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06673__A2 _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10665_ _05196_ _05198_ _05200_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12404_ _00905_ net456 u_cpu.rf_ram.memory\[116\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__I _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _05156_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A1 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12335_ _00836_ net364 u_cpu.rf_ram.memory\[120\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06425__A2 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05859__S1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__A3 _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12266_ _00767_ net355 u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10509__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09375__A1 _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08178__A2 _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11217_ _05557_ _05552_ _05559_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__S0 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12197_ _00711_ net298 u_cpu.rf_ram.memory\[127\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _05468_ _05514_ _05516_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__A1 _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11079_ u_cpu.rf_ram.memory\[83\]\[0\] _05471_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__I _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07689__A1 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout367_I net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08350__A2 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08438__I _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__I _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11237__A2 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout534_I net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02545_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08290_ u_cpu.rf_ram.memory\[29\]\[2\] _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06113__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07241_ _02749_ u_scanchain_local.module_data_in\[58\] _02788_ u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06664__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05797__I u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07172_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _02745_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08173__I _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__A1 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06123_ _01506_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11677__CLK net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07613__A1 u_cpu.rf_ram.memory\[78\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A2 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01698_ _01701_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08901__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout304 net305 net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout315 net320 net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11173__A1 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout326 net332 net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _04531_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout337 net338 net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout348 net352 net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06275__S1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05927__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10920__A1 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout359 net360 net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09118__A1 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09744_ u_cpu.rf_ram.memory\[33\]\[5\] _04475_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06956_ _02585_ u_cpu.rf_ram.rdata\[3\] _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05907_ _01555_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11476__A2 _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09675_ _04164_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06887_ _02460_ _02525_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12302__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A2 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08626_ _03638_ _03758_ _03765_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05838_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08348__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11228__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08557_ _02961_ _03595_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ _03020_ _03015_ _03022_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ _03346_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10987__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09841__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06655__A2 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07439_ _02932_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07852__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _05066_
+ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08083__I _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10739__A1 _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ _02914_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11400__A2 _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ u_cpu.rf_ram.memory\[32\]\[2\] _05027_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09907__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12120_ _00634_ net274 u_cpu.rf_ram.memory\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09357__A1 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12051_ _00565_ net15 u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11164__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11002_ u_cpu.rf_ram.memory\[79\]\[2\] _05424_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07907__A2 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06266__S1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10911__A1 _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09642__I _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11467__A2 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12953_ u_cpu.rf_ram_if.wdata1_r\[5\] net335 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11904_ _00426_ net271 u_cpu.rf_ram.memory\[60\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12884_ _01381_ net505 u_cpu.rf_ram.memory\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11219__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11835_ _00357_ net105 u_cpu.rf_ram.memory\[67\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06894__A2 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11766_ _00288_ net345 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10978__A1 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09832__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__C _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06646__A2 _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07843__A1 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10717_ _04679_ _04664_ _04791_ _04762_ _05242_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__06497__I2 u_cpu.rf_ram.memory\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11697_ _00219_ net452 u_cpu.rf_ram.memory\[43\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12945__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10648_ _04070_ _05184_ _05189_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10028__I _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout115_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _05109_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12318_ _00819_ net467 u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09348__A1 u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12249_ _00750_ net348 u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11155__A1 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09899__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06257__S1 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout484_I net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__A1 _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06810_ u_cpu.rf_ram.memory\[132\]\[7\] u_cpu.rf_ram.memory\[133\]\[7\] u_cpu.rf_ram.memory\[134\]\[7\]
+ u_cpu.rf_ram.memory\[135\]\[7\] _02101_ _01749_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06421__I2 u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ _03068_ _03168_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06741_ _02011_ _02382_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11458__A2 _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11734__D _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09520__A1 _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ u_cpu.rf_ram.memory\[92\]\[2\] _04301_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06672_ u_cpu.rf_ram.memory\[56\]\[6\] u_cpu.rf_ram.memory\[57\]\[6\] u_cpu.rf_ram.memory\[58\]\[6\]
+ u_cpu.rf_ram.memory\[59\]\[6\] _01652_ _01552_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12475__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08411_ _03581_ _03610_ _03619_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06724__I3 u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09391_ _04160_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_91_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _03346_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout28_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07834__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06637__A2 _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ u_cpu.rf_ram.memory\[64\]\[4\] _03530_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11322__I _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06193__S0 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__C _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07224_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_34_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07155_ _02714_ _02733_ _02734_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10441__I0 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06106_ u_cpu.rf_ram.memory\[140\]\[0\] u_cpu.rf_ram.memory\[141\]\[0\] u_cpu.rf_ram.memory\[142\]\[0\]
+ u_cpu.rf_ram.memory\[143\]\[0\] _01753_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07086_ _02680_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07601__A4 _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__A1 u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06037_ u_cpu.rf_ram.memory\[116\]\[0\] u_cpu.rf_ram.memory\[117\]\[0\] u_cpu.rf_ram.memory\[118\]\[0\]
+ u_cpu.rf_ram.memory\[119\]\[0\] _01684_ _01685_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout101 net103 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout112 net114 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout123 net142 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08011__A1 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout134 net135 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout145 net150 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout156 net157 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout167 net169 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08562__A2 _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout178 net179 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout189 net190 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07988_ _03349_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _04442_ _04460_ _04468_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06939_ _02575_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__A1 _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09658_ _04348_ _04415_ _04423_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08609_ _02949_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06876__A2 _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _04339_ _04377_ _04382_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11620_ _00142_ net437 u_cpu.rf_ram.memory\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__A1 u_cpu.rf_ram.memory\[77\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09814__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11551_ _03630_ _05766_ _05771_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07825__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ u_cpu.rf_ram.memory\[30\]\[2\] _05099_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11992__CLK net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11482_ _02890_ _05455_ _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10433_ _05057_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10188__A2 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _04970_ _05012_ _05014_ _05015_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08250__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12103_ _00617_ net264 u_cpu.rf_ram.memory\[137\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12348__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06800__A2 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10295_ _04951_ _04948_ _04953_ _04738_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12034_ _00548_ net419 u_cpu.rf_ram.memory\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06061__I _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08002__A1 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09750__A1 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12498__CLK net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10360__A2 _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12936_ u_cpu.rf_ram_if.wdata0_r\[1\] net340 u_cpu.rf_ram_if.wdata0_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12867_ _01364_ net500 u_cpu.rf_ram.memory\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06411__S1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06867__A2 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11818_ _00340_ net35 u_cpu.rf_ram.memory\[75\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12798_ _01295_ net412 u_cpu.rf_ram.memory\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06619__A2 _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07816__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _00271_ net429 u_cpu.rf_ram.memory\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout232_I net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09569__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11376__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10423__I0 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09547__I _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08241__A1 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08792__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _03969_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11715__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07911_ _01753_ _03296_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08891_ _03735_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07842_ u_cpu.rf_ram.memory\[50\]\[0\] _03246_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10351__A2 _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ _03129_ _03199_ _03201_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11865__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09512_ _04151_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06724_ u_cpu.rf_ram.memory\[136\]\[6\] u_cpu.rf_ram.memory\[137\]\[6\] u_cpu.rf_ram.memory\[138\]\[6\]
+ u_cpu.rf_ram.memory\[139\]\[6\] _01542_ _01544_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06158__I1 u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _04286_ _04287_ _04289_ _02563_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06655_ _01528_ _02297_ _01902_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06402__S1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09374_ _04241_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06586_ u_cpu.rf_ram.memory\[52\]\[5\] u_cpu.rf_ram.memory\[53\]\[5\] u_cpu.rf_ram.memory\[54\]\[5\]
+ u_cpu.rf_ram.memory\[55\]\[5\] _01647_ _02040_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07530__I _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08325_ _03564_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07807__A1 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ _03507_ _03515_ _03522_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ _02721_ u_scanchain_local.module_data_in\[53\] _02722_ u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ _03422_ _03470_ _03477_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05985__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07138_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _02719_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08783__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ _02664_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10590__A2 _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _04747_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08535__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__I1 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__I _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12790__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08299__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10982_ _05211_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12721_ _01218_ net155 u_cpu.rf_ram.memory\[99\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06849__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06765__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12652_ _01149_ net159 u_cpu.rf_ram.memory\[96\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12020__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11603_ _00125_ net416 u_cpu.rf_ram.memory\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12583_ _01081_ net327 u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11534_ u_cpu.rf_ram.memory\[89\]\[4\] _05758_ _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06056__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11465_ u_cpu.rf_ram.memory\[0\]\[0\] _05719_ _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05895__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09367__I u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10416_ _05047_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07026__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11396_ u_cpu.rf_ram.memory\[27\]\[5\] _05674_ _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10030__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10347_ _04908_ _04823_ _04999_ _04625_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06785__A1 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10278_ _04608_ _04714_ _04616_ _04835_ _04850_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11888__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09723__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12017_ _00531_ net61 u_cpu.rf_ram.memory\[141\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10242__S _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11530__A1 u_cpu.rf_ram.memory\[89\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__A2 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout182_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__S1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10097__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10976__I _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12919_ _01416_ net382 u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout447_I net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06440_ _02082_ _02084_ _02085_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08446__I _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07350__I _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06371_ u_cpu.rf_ram.memory\[8\]\[3\] u_cpu.rf_ram.memory\[9\]\[3\] u_cpu.rf_ram.memory\[10\]\[3\]
+ u_cpu.rf_ram.memory\[11\]\[3\] _02016_ _01564_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12513__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08110_ _03428_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09090_ u_cpu.rf_ram.memory\[130\]\[2\] _04055_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08462__A1 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ _03383_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10417__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__I _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08214__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10021__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09962__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ _04680_ _04681_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06776__A1 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10572__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08943_ u_cpu.rf_ram.memory\[49\]\[3\] _03962_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09714__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08517__A2 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ _03850_ _03914_ _03919_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06528__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11521__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10324__A2 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07825_ _03215_ _03233_ _03236_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09190__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06623__S1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _03139_ _03185_ _03190_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06707_ _02082_ _02349_ _02085_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10886__I _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07687_ _02933_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06585__B _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__I0 u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ u_cpu.rf_ram.memory\[90\]\[6\] _04271_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10883__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06638_ u_cpu.rf_ram.memory\[132\]\[5\] u_cpu.rf_ram.memory\[133\]\[5\] u_cpu.rf_ram.memory\[134\]\[5\]
+ u_cpu.rf_ram.memory\[135\]\[5\] _01993_ _02106_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09357_ _04228_ _03281_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12193__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06569_ _01547_ _02212_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06139__S0 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ u_cpu.rf_ram.memory\[63\]\[1\] _03553_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08453__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09288_ u_cpu.rf_ram.memory\[123\]\[4\] _04185_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08239_ u_cpu.rf_ram.memory\[66\]\[7\] _03494_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11250_ _05566_ _05572_ _05580_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07008__A2 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ _04861_ _04864_ _04867_ _04868_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08756__A2 _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _05484_ _05527_ _05535_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10132_ _04164_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09705__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08508__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _04629_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11512__A1 u_cpu.rf_ram.memory\[100\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06614__S1 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__I1 u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10079__A1 _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10796__I _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10965_ _05328_ _05389_ _05398_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12536__CLK net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12704_ _01201_ net154 u_cpu.rf_ram.memory\[103\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10896_ _05320_ _05351_ _05357_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12635_ _01132_ net152 u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A1 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12566_ _01064_ net310 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12686__CLK net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10251__A1 _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11517_ _03640_ _05743_ _05750_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12497_ _00998_ net492 u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06550__S0 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11448_ _05623_ _05706_ _05709_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08747__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11379_ _04861_ _05667_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09825__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10480__B _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout397_I net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05940_ _01511_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10306__A2 _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A2 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05871_ _01483_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07610_ _03088_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07722__A3 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08590_ _03731_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06930__A1 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07541_ u_cpu.rf_ram.memory\[1\]\[4\] _03043_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07472_ _02982_ _02988_ _02997_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08683__A1 _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07080__I _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09211_ u_cpu.rf_ram.memory\[126\]\[4\] _04132_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06423_ _01635_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10490__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09142_ u_cpu.rf_ram.memory\[22\]\[2\] _04091_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout10_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ u_cpu.rf_ram.memory\[24\]\[3\] u_cpu.rf_ram.memory\[25\]\[3\] u_cpu.rf_ram.memory\[26\]\[3\]
+ u_cpu.rf_ram.memory\[27\]\[3\] _01516_ _01774_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08904__I _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06297__I0 u_cpu.rf_ram.memory\[104\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _04003_ _04039_ _04045_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06285_ _01795_ _01918_ _01931_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_15_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10793__A2 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ u_cpu.rf_ram.memory\[129\]\[1\] _03373_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__A1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08738__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09975_ _04654_ _04666_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08926_ _03937_ _03946_ _03953_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06299__C _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09163__A2 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ u_cpu.rf_ram.memory\[14\]\[4\] _03906_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07174__A1 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12559__CLK net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _02939_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ u_cpu.rf_ram.memory\[71\]\[1\] _03865_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07739_ _03146_ _03171_ _03178_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10750_ _05215_ _05260_ _05267_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08086__I _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08674__A1 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09409_ _04264_ _04249_ _04265_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10681_ u_cpu.rf_ram.memory\[93\]\[4\] _05206_ _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06780__S0 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12420_ _00921_ net235 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06288__I0 u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12351_ _00852_ net364 u_cpu.rf_ram.memory\[121\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11240__I _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06532__S0 _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__A2 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ _05557_ _05607_ _05612_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12282_ _00783_ net398 u_cpu.rf_ram.memory\[91\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08729__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11233_ _03082_ _05455_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09926__A1 _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10536__A2 _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11164_ _03167_ _03197_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10115_ _04795_ _04796_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11095_ u_cpu.rf_ram.memory\[83\]\[5\] _05476_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10046_ _04706_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07165__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11997_ _00002_ net295 u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10948_ _05387_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08665__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout145_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10879_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _05341_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06140__A2 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12618_ _01115_ net146 u_cpu.rf_ram.memory\[93\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08968__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12549_ _01049_ net173 u_cpu.rf_ram.memory\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout312_I net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__S0 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A1 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10775__A2 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06244__I _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06070_ _01704_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07640__A2 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09393__A2 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout508 net509 net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout519 net523 net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09760_ _04491_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06972_ _01496_ _02586_ _02601_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ _03752_ _03808_ _03816_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05923_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09691_ _04446_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08642_ u_cpu.rf_ram.memory\[15\]\[2\] _03775_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05854_ _01502_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10430__S _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12851__CLK net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08573_ u_cpu.rf_ram.memory\[53\]\[6\] _03722_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05785_ _01436_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _01437_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_82_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07524_ u_cpu.cpu.immdec.imm11_7\[2\] _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06419__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07455_ _02986_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06406_ _01568_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08634__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08408__A1 u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07386_ _02902_ u_cpu.rf_ram_if.wdata0_r\[4\] _02930_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_52_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ _02945_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10215__A1 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06337_ _01958_ _01970_ _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09081__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10766__A2 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09056_ u_cpu.rf_ram.memory\[132\]\[5\] _04031_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12231__CLK net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06268_ _01537_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07631__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ u_cpu.rf_ram.memory\[119\]\[3\] _03362_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06199_ _01618_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05993__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06037__I3 u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06198__A2 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__A2 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12381__CLK net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09958_ _04609_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08909_ _03941_ _03928_ _03942_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09889_ u_cpu.rf_ram.memory\[113\]\[1\] _04586_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _00442_ net220 u_cpu.rf_ram.memory\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__A2 _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06757__C _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11851_ _00373_ net105 u_cpu.rf_ram.memory\[65\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11235__I _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10802_ _05294_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08647__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11782_ _00304_ net269 u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10733_ u_cpu.cpu.immdec.imm30_25\[0\] _04670_ _05224_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06753__S0 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10664_ u_cpu.rf_ram.memory\[93\]\[0\] _05199_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08544__I _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07870__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06492__C _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12403_ _00904_ net455 u_cpu.rf_ram.memory\[116\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10206__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09072__A1 u_cpu.rf_ram.memory\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _05107_ _05110_ _05155_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06064__I _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12334_ _00835_ net364 u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06681__I0 u_cpu.rf_ram.memory\[100\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06999__I _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12265_ _00766_ net358 u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12724__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07096__S _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11216_ u_cpu.rf_ram.memory\[85\]\[2\] _05558_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09375__A2 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06808__S1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12196_ _00710_ net296 u_cpu.rf_ram.memory\[127\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07386__A1 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11182__A2 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11147_ u_cpu.rf_ram.memory\[84\]\[0\] _05515_ _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09127__A2 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12874__CLK net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11078_ _05469_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07138__A1 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10029_ _04686_ _04714_ _04620_ _04716_ _04717_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07689__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__A1 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout262_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__I3 u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12104__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11145__I _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10189__C _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__A1 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09835__B1 _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout527_I net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06744__S0 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ _02696_ _02804_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12254__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07171_ _02745_ _02746_ _02747_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10748__A2 _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06122_ _01497_ _01645_ _01770_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07613__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06053_ _01484_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07377__A1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout305 net306 net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout316 net318 net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11173__A2 _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06424__I0 u_cpu.rf_ram.memory\[116\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _04532_ _04535_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout327 net331 net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout338 net342 net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout349 net352 net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05927__A2 _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09743_ _04438_ _04471_ _04478_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06955_ _02584_ _02589_ _02590_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05906_ _01532_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09674_ _04433_ _04428_ _04435_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06886_ _02517_ _02521_ _02523_ _02524_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08877__A1 u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ u_cpu.rf_ram.memory\[9\]\[4\] _03762_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05837_ _01486_ _01487_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08629__A1 u_cpu.rf_ram.memory\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06149__I _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08556_ _03679_ _03707_ _03716_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07507_ u_cpu.rf_ram.memory\[20\]\[2\] _03021_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _03673_ _03663_ _03674_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07301__A1 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06735__S0 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05988__I _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10987__A2 _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07438_ _02974_ _02966_ _02975_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07852__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11621__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _02901_ _02915_ _02916_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10739__A2 _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09108_ _04062_ _04065_ _04067_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _05022_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08801__A1 u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06663__I0 u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09039_ _04009_ _04016_ _04024_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09357__A2 _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12050_ _00564_ net36 u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11771__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07368__A1 u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11001_ _05419_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06415__I0 u_cpu.rf_ram.memory\[124\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06591__A2 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12952_ u_cpu.rf_ram_if.wdata1_r\[4\] net341 u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08539__I _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08868__A1 u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11903_ _00425_ net90 u_cpu.rf_ram.memory\[60\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12883_ _01380_ net505 u_cpu.rf_ram.memory\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07540__A1 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12001__D _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12277__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11834_ _00356_ net19 u_cpu.rf_ram.memory\[68\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11765_ _00287_ net301 u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09293__A1 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05898__I _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06726__S0 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10716_ _04722_ _04902_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11696_ _00218_ net452 u_cpu.rf_ram.memory\[43\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07843__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10647_ u_cpu.rf_ram.memory\[2\]\[2\] _05188_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10578_ _05145_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12317_ _00818_ net487 u_cpu.rf_ram.memory\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__A2 _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12248_ _00749_ net348 u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12179_ _00693_ net185 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10979__I _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06740_ u_cpu.rf_ram.memory\[4\]\[7\] u_cpu.rf_ram.memory\[5\]\[7\] u_cpu.rf_ram.memory\[6\]\[7\]
+ u_cpu.rf_ram.memory\[7\]\[7\] _01561_ _01564_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__A1 u_cpu.rf_ram.memory\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07353__I _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06671_ _01919_ _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ u_cpu.rf_ram.memory\[19\]\[7\] _03608_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _04251_ _04248_ _04252_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08341_ _03575_ _03565_ _03576_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11644__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08272_ _03503_ _03526_ _03532_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07834__A2 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06193__S1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05845__A1 _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07223_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_69_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11794__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _02721_ u_scanchain_local.module_data_in\[43\] _02722_ u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11394__A2 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06105_ _01748_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07085_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_dbus_dat\[23\] _02677_ _02680_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07528__I _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06270__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09944__S _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06036_ _01637_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout102 net103 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08011__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout135 net140 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout146 net149 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06022__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout157 net158 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07070__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout168 net169 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout179 net180 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07987_ _02944_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09726_ u_cpu.rf_ram.memory\[116\]\[6\] _04463_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06938_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _02513_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10657__A1 u_cpu.rf_ram.memory\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09657_ u_cpu.rf_ram.memory\[112\]\[6\] _04418_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06869_ _02504_ _02501_ _02506_ _02508_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_55_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03752_ _03733_ _03753_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09588_ u_cpu.rf_ram.memory\[121\]\[2\] _04381_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _03705_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11550_ u_cpu.rf_ram.memory\[23\]\[2\] _05770_ _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11082__A1 u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07825__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _05094_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11481_ _02982_ _05719_ _05728_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10129__I _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _05054_
+ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07589__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11385__A2 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__I0 u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ u_cpu.cpu.immdec.imm19_12_20\[8\] _04947_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08250__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12102_ _00616_ net261 u_cpu.rf_ram.memory\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06261__A1 _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10294_ u_cpu.cpu.immdec.imm19_12_20\[2\] _04949_ _04952_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12033_ _00547_ net419 u_cpu.rf_ram.memory\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08002__A2 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07061__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10896__A1 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09750__A2 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07761__A1 u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10648__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09502__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12935_ _01431_ net314 u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06167__I2 u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10112__A3 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12912__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12866_ _01363_ net501 u_cpu.rf_ram.memory\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A2 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11817_ _00339_ net35 u_cpu.rf_ram.memory\[75\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09266__A1 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11423__I _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12797_ _01294_ net412 u_cpu.rf_ram.memory\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11073__A1 u_cpu.rf_ram.memory\[107\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11748_ _00270_ net432 u_cpu.rf_ram.memory\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07816__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11679_ _00201_ net391 u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09828__I _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09569__A2 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08241__A2 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10584__B1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06252__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11128__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07910_ _02886_ _03295_ _03296_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08890_ _03925_ _03927_ _03929_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07841_ _03244_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12442__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__A2 _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__A1 u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07772_ u_cpu.rf_ram.memory\[43\]\[0\] _03200_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08179__I _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10639__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09511_ _04264_ _04322_ _04331_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06723_ _01763_ _02365_ _01485_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07504__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06158__I2 u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12592__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09442_ _04288_ _02548_ _02495_ _02487_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06654_ u_cpu.rf_ram.memory\[0\]\[6\] u_cpu.rf_ram.memory\[1\]\[6\] u_cpu.rf_ram.memory\[2\]\[6\]
+ u_cpu.rf_ram.memory\[3\]\[6\] _01529_ _01900_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout40_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08907__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07811__I _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ _03270_ _04228_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09257__A1 u_cpu.rf_ram.memory\[124\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06585_ _01651_ _02228_ _01520_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11064__A1 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08324_ _03082_ _03168_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07807__A2 _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ u_cpu.rf_ram.memory\[65\]\[5\] _03518_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08480__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07206_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _02775_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06491__A1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ u_cpu.rf_ram.memory\[68\]\[5\] _03473_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ _02715_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _02710_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07068_ _02670_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09980__A2 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11119__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06019_ _01616_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09473__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07743__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12935__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08089__I _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _04444_ _04448_ _04457_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10981_ _05409_ _05401_ _05410_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09496__A1 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08299__A2 _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12720_ _01217_ net156 u_cpu.rf_ram.memory\[99\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12651_ _01148_ net195 u_cpu.rf_ram.memory\[96\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__A1 u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11602_ _00124_ net416 u_cpu.rf_ram.memory\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11055__A1 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12582_ _01080_ net327 u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05809__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11533_ _03634_ _05754_ _05760_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12315__CLK net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__B _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09648__I _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11464_ _05717_ _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10415_ _02530_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11395_ _05630_ _05670_ _05677_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06072__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10346_ _04749_ _04781_ _04765_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10030__A2 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07982__A1 _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10277_ _04931_ _04934_ _04937_ _04686_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12016_ _00530_ net57 u_cpu.rf_ram.memory\[141\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06537__A2 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11530__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout175_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09487__A1 _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10097__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12918_ _01415_ net382 u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout342_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12849_ _01346_ net436 u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11046__A1 u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06370_ _01503_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10254__C1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08040_ _03383_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__A2 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__A1 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10021__A2 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09962__A2 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09991_ _04619_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06776__A2 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11832__CLK net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12958__CLK net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08942_ _03932_ _03958_ _03963_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout88_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08873_ u_cpu.rf_ram.memory\[138\]\[2\] _03918_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06528__A2 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06084__S0 _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07824_ u_cpu.rf_ram.memory\[47\]\[1\] _03234_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11982__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09478__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07755_ u_cpu.rf_ram.memory\[41\]\[2\] _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06706_ u_cpu.rf_ram.memory\[84\]\[6\] u_cpu.rf_ram.memory\[85\]\[6\] u_cpu.rf_ram.memory\[86\]\[6\]
+ u_cpu.rf_ram.memory\[87\]\[6\] _01684_ _02083_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07686_ _03142_ _03134_ _03143_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09425_ _04260_ _04268_ _04275_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06637_ _01539_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11037__A1 u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06157__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06568_ u_cpu.rf_ram.memory\[8\]\[5\] u_cpu.rf_ram.memory\[9\]\[5\] u_cpu.rf_ram.memory\[10\]\[5\]
+ u_cpu.rf_ram.memory\[11\]\[5\] _02016_ _01507_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09356_ _02505_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06139__S1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08307_ _03493_ _03552_ _03554_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _04165_ _04181_ _04187_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09650__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06499_ u_cpu.rf_ram.memory\[48\]\[4\] u_cpu.rf_ram.memory\[49\]\[4\] u_cpu.rf_ram.memory\[50\]\[4\]
+ u_cpu.rf_ram.memory\[51\]\[4\] _01636_ _01927_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06303__I2 u_cpu.rf_ram.memory\[122\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _03352_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12488__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ _02946_ _03458_ _03466_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09402__A1 u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08205__A2 _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10548__B1 _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _04686_ _04722_ _04684_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11180_ u_cpu.rf_ram.memory\[59\]\[6\] _05530_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__A2 _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07964__A1 u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _04807_ _04802_ _04809_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09705__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _04747_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_62_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07716__A1 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11512__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09469__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06776__B _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11276__A1 u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10079__A2 _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10964_ u_cpu.rf_ram.memory\[104\]\[7\] _05387_ _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12703_ _01200_ net154 u_cpu.rf_ram.memory\[103\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10895_ u_cpu.rf_ram.memory\[101\]\[3\] _05355_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08692__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12634_ _01131_ net151 u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11705__CLK net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__A1 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12565_ _01063_ net309 u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11516_ u_cpu.rf_ram.memory\[100\]\[5\] _05746_ _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10251__A2 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12496_ _00997_ net492 u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06550__S1 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11447_ u_cpu.rf_ram.memory\[24\]\[1\] _05707_ _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11200__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10003__A2 _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11378_ u_cpu.cpu.ctrl.i_iscomp _04601_ _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10329_ u_cpu.cpu.immdec.imm19_12_20\[6\] _04698_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout292_I net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07707__A1 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10306__A3 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ u_cpu.rf_ram.memory\[24\]\[0\] u_cpu.rf_ram.memory\[25\]\[0\] u_cpu.rf_ram.memory\[26\]\[0\]
+ u_cpu.rf_ram.memory\[27\]\[0\] _01516_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08380__A1 u_cpu.rf_ram.memory\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07722__A4 _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ _02928_ _03039_ _03045_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07471_ u_cpu.rf_ram.memory\[81\]\[7\] _02986_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09880__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__A2 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06422_ _02065_ _02067_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09210_ _04093_ _04128_ _04134_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10490__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12630__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ _04084_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06353_ _01500_ _01998_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10428__S _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08435__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09632__A1 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09072_ u_cpu.rf_ram.memory\[131\]\[3\] _04043_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08192__I _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06284_ _01921_ _01923_ _01925_ _01930_ _01642_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08023_ _03326_ _03372_ _03374_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12780__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08199__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09935__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07946__A1 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09974_ _04655_ _04665_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07536__I _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12010__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09952__S _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08925_ u_cpu.rf_ram.memory\[137\]\[4\] _03950_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__A1 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03635_ _03902_ _03908_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _03222_ _03212_ _03223_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05999_ _01600_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08787_ _03843_ _03864_ _03866_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12160__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__B _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07738_ u_cpu.rf_ram.memory\[51\]\[5\] _03174_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08123__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07669_ _03103_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08674__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ u_cpu.rf_ram.memory\[91\]\[7\] _04247_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10680_ _05211_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__S1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09339_ u_cpu.rf_ram.memory\[36\]\[0\] _04218_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11878__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12350_ _00851_ net361 u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11301_ u_cpu.rf_ram.memory\[87\]\[2\] _05611_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06532__S1 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12281_ _00782_ net380 u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11232_ _05568_ _05553_ _05569_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09926__A2 _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__A1 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11163_ _05486_ _05515_ _05524_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10114_ _04700_ _04779_ _04679_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11094_ _05214_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11497__A1 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07890__B _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10045_ _04731_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__I _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08362__A1 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06599__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11249__A1 u_cpu.rf_ram.memory\[110\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__I0 u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11996_ _00001_ net295 u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08114__A1 _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12653__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10947_ _05387_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09862__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08665__A2 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09862__B2 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06220__S0 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10878_ _05346_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06771__S1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12617_ _01114_ net152 u_cpu.rf_ram.memory\[93\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09614__A1 u_cpu.rf_ram.memory\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13009__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout138_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06428__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__A1 _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12548_ _01048_ net172 u_cpu.rf_ram.memory\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__A2 _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06523__S1 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A2 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout305_I net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12479_ _00980_ net240 u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12033__CLK net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07928__A1 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout509 net510 net509 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06600__A1 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06971_ u_cpu.rf_ram_if.rdata0\[2\] _02599_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08710_ u_cpu.rf_ram.memory\[140\]\[6\] _03811_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11488__A1 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05922_ _01505_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09690_ _03166_ _04426_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08641_ _03770_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05853_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05784_ u_cpu.rf_ram_if.rcnt\[0\] _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08572_ _03675_ _03719_ _03726_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07523_ _03031_ _03016_ _03032_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09853__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09853__B2 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06506__I2 u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07454_ _02986_ _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06405_ _01937_ _02050_ _01654_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _02903_ u_cpu.rf_ram_if.wdata1_r\[4\] _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09605__A1 u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08408__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09124_ _04077_ _04066_ _04078_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06336_ _01974_ _01976_ _01978_ _01981_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__10215__A2 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09081__A2 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _04005_ _04027_ _04034_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06267_ _01599_ _01913_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08006_ _03337_ _03358_ _03363_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06198_ _01494_ _01833_ _01845_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12526__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06198__A3 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08592__A1 _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09957_ _04646_ _04648_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ u_cpu.rf_ram.memory\[39\]\[6\] _03933_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09888_ _04425_ _04585_ _04587_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08344__A1 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08839_ _03857_ _03890_ _03897_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10151__A1 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11850_ _00372_ net106 u_cpu.rf_ram.memory\[66\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05953__I0 u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10801_ _05202_ _05295_ _05298_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08647__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11781_ _00303_ net273 u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06202__S0 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10732_ _04720_ _04862_ _05255_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06753__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10663_ _05197_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12402_ _00903_ net455 u_cpu.rf_ram.memory\[116\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12056__CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10206__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06345__I _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10594_ _01454_ _05153_ _05154_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09072__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12333_ _00834_ net479 u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06830__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06681__I1 u_cpu.rf_ram.memory\[101\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12264_ _00765_ net355 u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11215_ _05551_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12195_ _00709_ net293 u_cpu.rf_ram.memory\[127\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08583__A1 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ _05513_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10390__A1 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11077_ _05469_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08335__A1 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10028_ _04598_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10142__A1 u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08886__A2 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06897__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10693__A2 _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout255_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11979_ _00501_ net221 u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09835__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09835__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06744__S1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout422_I net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06255__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07170_ _02684_ u_scanchain_local.module_data_in\[46\] _02730_ u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ _01744_ _01769_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06052_ u_cpu.rf_ram.memory\[88\]\[0\] u_cpu.rf_ram.memory\[89\]\[0\] u_cpu.rf_ram.memory\[90\]\[0\]
+ u_cpu.rf_ram.memory\[91\]\[0\] _01699_ _01700_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07377__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout306 net371 net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08574__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ u_arbiter.i_wb_cpu_rdt\[8\] _04533_ _04534_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xfanout317 net318 net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout328 net331 net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout339 net342 net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ u_cpu.rf_ram.memory\[33\]\[4\] _04475_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10441__S _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout70_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06954_ _02587_ u_cpu.rf_ram_if.rdata1\[2\] _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07814__I _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05905_ u_cpu.rf_ram.memory\[0\]\[0\] u_cpu.rf_ram.memory\[1\]\[0\] u_cpu.rf_ram.memory\[2\]\[0\]
+ u_cpu.rf_ram.memory\[3\]\[0\] _01550_ _01553_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10133__A1 u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09673_ u_cpu.rf_ram.memory\[122\]\[2\] _04434_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06885_ _01443_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08877__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _03635_ _03758_ _03764_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06432__S0 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05836_ u_cpu.cpu.immdec.imm24_20\[2\] _01473_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08555_ u_cpu.rf_ram.memory\[54\]\[7\] _03705_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08629__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09826__A1 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12079__CLK net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07506_ _03014_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ u_cpu.rf_ram.memory\[57\]\[4\] _03669_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06735__S1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07437_ u_cpu.rf_ram.memory\[21\]\[3\] _02972_ _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ u_cpu.rf_ram.memory\[82\]\[1\] _02909_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09054__A2 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09107_ u_cpu.rf_ram.memory\[12\]\[0\] _04066_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06319_ u_cpu.rf_ram.memory\[80\]\[2\] u_cpu.rf_ram.memory\[81\]\[2\] u_cpu.rf_ram.memory\[82\]\[2\]
+ u_cpu.rf_ram.memory\[83\]\[2\] _01706_ _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07299_ _02558_ u_cpu.cpu.decode.opcode\[1\] _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06112__I0 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08801__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09038_ u_cpu.rf_ram.memory\[133\]\[6\] _04019_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11916__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10415__I _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07368__A2 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11000_ _05404_ _05420_ _05423_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08317__A1 u_cpu.rf_ram.memory\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06591__A3 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12951_ u_cpu.rf_ram_if.wdata1_r\[3\] net341 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__A1 _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08868__A2 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10150__I _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11902_ _00424_ net90 u_cpu.rf_ram.memory\[60\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12882_ _01379_ net502 u_cpu.rf_ram.memory\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11833_ _00355_ net12 u_cpu.rf_ram.memory\[68\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09817__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09817__B2 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _00286_ net300 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06726__S1 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10715_ _05239_ _05240_ _04964_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11695_ _00217_ net402 u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06075__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10646_ _05183_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09045__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10577_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _05144_ _05139_ u_cpu.cpu.ctrl.o_ibus_adr\[25\]
+ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11596__CLK net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12316_ _00817_ net465 u_cpu.rf_ram.memory\[35\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12841__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12247_ _00748_ net361 u_cpu.rf_ram.memory\[123\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08556__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12178_ _00692_ net424 u_cpu.rf_ram.memory\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11357__S _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11129_ _05473_ _05501_ _05504_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12991__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A1 u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout372_I net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06670_ u_cpu.rf_ram.memory\[60\]\[6\] u_cpu.rf_ram.memory\[61\]\[6\] u_cpu.rf_ram.memory\[62\]\[6\]
+ u_cpu.rf_ram.memory\[63\]\[6\] _01668_ _02034_ _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12221__CLK net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10995__I _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09808__A1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08340_ u_cpu.rf_ram.memory\[62\]\[4\] _03571_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ u_cpu.rf_ram.memory\[64\]\[3\] _03530_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07295__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07222_ _02724_ _02787_ _02789_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09036__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _02732_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10436__S _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01541_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08795__A1 u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07084_ _02679_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06035_ _01635_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_86_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__A1 u_cpu.rf_ram.memory\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout103 net104 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout114 net117 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout125 net126 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout136 net139 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout147 net149 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout158 net160 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06022__A2 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07070__I1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _03347_ _03331_ _03348_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout169 net180 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09725_ _04440_ _04460_ _04467_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06937_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _02500_ _02574_ _02575_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__10106__A1 _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10657__A2 _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _04346_ _04415_ _04422_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06868_ _02460_ _02507_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08607_ u_cpu.rf_ram.memory\[52\]\[6\] _03740_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05819_ u_cpu.rf_ram_if.rtrig0 _01455_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09587_ _04376_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06799_ u_cpu.rf_ram.memory\[68\]\[7\] u_cpu.rf_ram.memory\[69\]\[7\] u_cpu.rf_ram.memory\[70\]\[7\]
+ u_cpu.rf_ram.memory\[71\]\[7\] _01712_ _01713_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12714__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05999__I _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10409__A2 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08538_ _03705_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07286__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06333__I0 u_cpu.rf_ram.memory\[76\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _03325_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10500_ _04805_ _05095_ _05098_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11480_ u_cpu.rf_ram.memory\[0\]\[7\] _05717_ _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12864__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _05056_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05948__B _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07589__A2 _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__A1 u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10362_ _02617_ _02534_ _05013_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10593__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12101_ _00615_ net264 u_cpu.rf_ram.memory\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10293_ _04946_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12032_ _00546_ net419 u_cpu.rf_ram.memory\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10345__A1 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07061__I1 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10896__A2 _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12244__CLK net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10648__A2 _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12934_ _01430_ net378 u_cpu.rf_ram.memory\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12947__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12865_ _01362_ net501 u_cpu.rf_ram.memory\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12394__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11816_ _00338_ net35 u_cpu.rf_ram.memory\[75\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12796_ _01293_ net412 u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07277__A1 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11747_ _00269_ net432 u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11073__A2 _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11678_ _00200_ net391 u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__A1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout120_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10629_ u_cpu.rf_ram.memory\[3\]\[3\] _05176_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10256__S _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout218_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06627__I1 u_cpu.rf_ram.memory\[77\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06252__A2 _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10336__A1 _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07201__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07840_ _03244_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07771_ _03198_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11611__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12737__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09510_ u_cpu.rf_ram.memory\[34\]\[7\] _04320_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06722_ u_cpu.rf_ram.memory\[132\]\[6\] u_cpu.rf_ram.memory\[133\]\[6\] u_cpu.rf_ram.memory\[134\]\[6\]
+ u_cpu.rf_ram.memory\[135\]\[6\] _02101_ _01749_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10639__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07504__A2 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ u_cpu.cpu.alu.cmp_r _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06653_ _02011_ _02295_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__B _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09372_ _04239_ _03294_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08195__I _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09257__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06584_ u_cpu.rf_ram.memory\[56\]\[5\] u_cpu.rf_ram.memory\[57\]\[5\] u_cpu.rf_ram.memory\[58\]\[5\]
+ u_cpu.rf_ram.memory\[59\]\[5\] _01652_ _01812_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _03325_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11064__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__I0 u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10811__A2 _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08254_ _03505_ _03514_ _03521_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _02769_ _02765_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _03420_ _03469_ _03476_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07136_ _02714_ _02717_ _02718_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07440__A1 u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_dbus_dat\[15\] _02665_ _02670_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09754__I _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06018_ _01581_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07969_ _03334_ _03330_ _03335_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09708_ u_cpu.rf_ram.memory\[115\]\[7\] _04446_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10980_ u_cpu.rf_ram.memory\[99\]\[3\] _05407_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09496__A2 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ u_cpu.rf_ram.memory\[11\]\[7\] _04401_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _01147_ net195 u_cpu.rf_ram.memory\[96\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11601_ _00123_ net416 u_cpu.rf_ram.memory\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07259__A1 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11055__A2 _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12581_ _01079_ net327 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11532_ u_cpu.rf_ram.memory\[89\]\[3\] _05758_ _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05809__A2 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06482__A2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11463_ _05717_ _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10076__S _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08759__A1 u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10414_ _02869_ _04290_ _05046_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11394_ u_cpu.rf_ram.memory\[27\]\[4\] _05674_ _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07431__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _04908_ _04963_ _04617_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09664__I _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__A1 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10276_ _04623_ _04935_ _04936_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11634__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12015_ _00529_ net45 u_cpu.rf_ram.memory\[141\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07195__B1 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11784__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12917_ _01414_ net175 u_cpu.rf_ram.memory\[100\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout168_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12848_ _01345_ net435 u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06170__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout335_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12779_ _01276_ net18 u_cpu.rf_ram.memory\[69\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08998__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10254__C2 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__I3 u_cpu.rf_ram.memory\[95\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout502_I net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__A2 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07359__I _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__A1 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _03277_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ u_cpu.rf_ram.memory\[49\]\[2\] _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10309__A1 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05984__A1 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09175__A1 u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06608__S0 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ _03913_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08922__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ _03210_ _03233_ _03235_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06084__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07754_ _03184_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09478__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06705_ _01678_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07685_ u_cpu.rf_ram.memory\[45\]\[3\] _03140_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06536__I0 u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11344__I _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09424_ u_cpu.rf_ram.memory\[90\]\[5\] _04271_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06000__I2 u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06636_ u_cpu.rf_ram.memory\[128\]\[5\] u_cpu.rf_ram.memory\[129\]\[5\] u_cpu.rf_ram.memory\[130\]\[5\]
+ u_cpu.rf_ram.memory\[131\]\[5\] _01542_ _01544_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11037__A2 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04177_ _04218_ _04227_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06567_ _01785_ _02210_ _01902_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08306_ u_cpu.rf_ram.memory\[63\]\[0\] _03553_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08989__A1 u_cpu.rf_ram.memory\[135\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09286_ u_cpu.rf_ram.memory\[123\]\[3\] _04185_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06498_ _02039_ _02142_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09650__A2 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ _03509_ _03496_ _03510_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06464__A2 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ u_cpu.rf_ram.memory\[6\]\[6\] _03461_ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09402__A2 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10548__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11657__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07119_ _02702_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12902__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08099_ _03346_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10130_ u_cpu.rf_ram.memory\[114\]\[2\] _04808_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06767__A3 _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07964__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _04602_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06122__B _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__A1 _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10720__A1 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10963_ _05326_ _05389_ _05397_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10079__A3 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11254__I _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12702_ _01199_ net154 u_cpu.rf_ram.memory\[103\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10894_ _05317_ _05351_ _05356_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12633_ _01130_ net194 u_cpu.rf_ram.memory\[97\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11028__A2 _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__B _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12564_ _01062_ net309 u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12432__CLK net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10787__A1 u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09641__A2 _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _03637_ _05742_ _05749_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07652__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12495_ _00996_ net316 u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06083__I _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11446_ _05618_ _05706_ _05708_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11200__A2 _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12582__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11377_ _05665_ _05666_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10328_ _04620_ _04971_ _04982_ _04600_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11429__I _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09157__A1 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10259_ _04891_ _04749_ _04910_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09952__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10711__A1 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout285_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08380__A2 _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11267__A2 _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout452_I net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08132__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07470_ _02980_ _02988_ _02996_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06421_ u_cpu.rf_ram.memory\[112\]\[3\] u_cpu.rf_ram.memory\[113\]\[3\] u_cpu.rf_ram.memory\[114\]\[3\]
+ u_cpu.rf_ram.memory\[115\]\[3\] _02066_ _01840_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11019__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07891__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _03738_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06352_ u_cpu.rf_ram.memory\[28\]\[3\] u_cpu.rf_ram.memory\[29\]\[3\] u_cpu.rf_ram.memory\[30\]\[3\]
+ u_cpu.rf_ram.memory\[31\]\[3\] _01504_ _01771_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07643__A1 _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ _04000_ _04039_ _04044_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06283_ _01926_ _01928_ _01929_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06297__I2 u_cpu.rf_ram.memory\[106\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12925__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ u_cpu.rf_ram.memory\[129\]\[0\] _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__A1 u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08199__A2 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10250__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09973_ _04662_ _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__A1 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09148__A1 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08924_ _03935_ _03946_ _03952_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09699__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09943__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08855_ u_cpu.rf_ram.memory\[14\]\[3\] _03906_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12305__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07806_ u_cpu.rf_ram.memory\[48\]\[4\] _03218_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08786_ u_cpu.rf_ram.memory\[71\]\[0\] _03865_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _01568_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07552__I _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11258__A2 _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _03144_ _03170_ _03177_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09320__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08123__A2 _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _02907_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09871__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09407_ _04176_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06619_ _02082_ _02262_ _02085_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07599_ _03033_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_16_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09479__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09338_ _04216_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10769__A1 u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07634__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11430__A2 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06288__I2 u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ u_cpu.rf_ram.memory\[124\]\[6\] _04162_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11300_ _05606_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12280_ _00781_ net380 u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09387__A1 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11231_ u_cpu.rf_ram.memory\[85\]\[7\] _05551_ _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11194__A1 _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07937__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11162_ u_cpu.rf_ram.memory\[84\]\[7\] _05513_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05948__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10941__A1 _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09139__A1 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10113_ _04728_ _04794_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11093_ _05480_ _05470_ _05481_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10044_ _04708_ _04630_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08362__A2 _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11995_ _00000_ net291 u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09311__A1 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08114__A2 _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10946_ _03327_ _05374_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09862__A2 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06220__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10877_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _05341_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12948__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12616_ _01113_ net159 u_cpu.rf_ram.memory\[93\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12547_ _01047_ net187 u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06428__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11421__A2 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12478_ _00979_ net240 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11972__CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout200_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _05693_ _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08050__A1 _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05939__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10932__A1 _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__A2 _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10063__I _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06970_ _01496_ _02475_ _02600_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05921_ _01569_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06697__B _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07156__A3 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09550__A1 u_cpu.rf_ram.memory\[120\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ _03628_ _03771_ _03774_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05852_ u_cpu.raddr\[0\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__B2 _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07372__I _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12478__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ u_cpu.rf_ram.memory\[53\]\[5\] _03722_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09302__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07522_ u_cpu.rf_ram.memory\[20\]\[7\] _03014_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10999__A1 u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07453_ _02899_ _02985_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10439__S _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ u_cpu.rf_ram.memory\[96\]\[3\] u_cpu.rf_ram.memory\[97\]\[3\] u_cpu.rf_ram.memory\[98\]\[3\]
+ u_cpu.rf_ram.memory\[99\]\[3\] _01938_ _01824_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07384_ _02901_ _02928_ _02929_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09605__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09123_ u_cpu.rf_ram.memory\[12\]\[5\] _04071_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07616__A1 _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06335_ _01577_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10238__I _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ u_cpu.rf_ram.memory\[132\]\[4\] _04031_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06266_ u_cpu.rf_ram.memory\[40\]\[2\] u_cpu.rf_ram.memory\[41\]\[2\] u_cpu.rf_ram.memory\[42\]\[2\]
+ u_cpu.rf_ram.memory\[43\]\[2\] _01569_ _01601_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09369__A1 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ u_cpu.rf_ram.memory\[119\]\[2\] _03362_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06197_ _01835_ _01839_ _01842_ _01844_ _01689_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10923__A1 u_cpu.rf_ram.memory\[102\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08592__A2 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09956_ _03275_ u_arbiter.i_wb_cpu_rdt\[12\] _04647_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08907_ _03751_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__A2 _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09887_ u_cpu.rf_ram.memory\[113\]\[0\] _04586_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08344__A2 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08838_ u_cpu.rf_ram.memory\[143\]\[5\] _03893_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10151__A2 _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08769_ u_cpu.rf_ram.memory\[73\]\[3\] _03851_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05953__I1 u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11845__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10800_ u_cpu.rf_ram.memory\[96\]\[1\] _05296_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11780_ _00302_ net268 u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09844__A2 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10731_ _04740_ _04762_ _05254_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06202__S1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10662_ _05197_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09002__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12401_ _00902_ net455 u_cpu.rf_ram.memory\[116\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07607__A1 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10593_ _02477_ _02548_ _01454_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12332_ _00833_ net454 u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__A1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12263_ _00764_ net360 u_cpu.rf_ram.memory\[37\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06681__I2 u_cpu.rf_ram.memory\[102\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06361__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11214_ _05204_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08032__A1 _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06269__S1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12194_ _00708_ net268 u_cpu.rf_ram.memory\[128\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10914__A1 _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08583__A2 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ _05513_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06594__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09672__I _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12620__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11076_ _04295_ _03480_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A1 u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08335__A2 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10027_ _04596_ u_arbiter.i_wb_cpu_rdt\[5\] _04715_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06897__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12770__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11978_ _00500_ net67 u_cpu.rf_ram.memory\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09835__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout150_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ u_cpu.rf_ram.memory\[103\]\[0\] _05377_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout248_I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10486__C _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09599__A1 _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06120_ _01751_ _01757_ _01762_ _01767_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06051_ _01607_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12150__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06672__I2 u_cpu.rf_ram.memory\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07367__I _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11718__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08023__A1 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__A1 _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout307 net312 net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09810_ _04518_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09771__A1 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08574__A2 _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout318 net319 net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout329 net330 net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06585__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09582__I _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _04436_ _04471_ _04477_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06953_ _02585_ u_cpu.rf_ram.rdata\[2\] _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09523__A1 u_cpu.rf_ram.memory\[117\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ _01552_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09672_ _04427_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06337__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06884_ _02490_ _02522_ _02464_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11330__A1 u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08623_ u_cpu.rf_ram.memory\[9\]\[3\] _03762_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05835_ u_cpu.cpu.immdec.imm19_12_20\[6\] _01440_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06432__S1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _03677_ _03707_ _03715_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09826__A2 _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ _02920_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_23_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08485_ _03343_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07436_ _02926_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07367_ _02914_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11397__A1 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ _04064_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06318_ _01585_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08661__I _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ _02480_ u_cpu.cpu.bufreg.c_r _02850_ _02851_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06499__S1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09037_ _04007_ _04016_ _04023_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06249_ _01887_ _01889_ _01893_ _01895_ _01490_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A1 _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09762__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A1 _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _04613_ _04630_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__A2 _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12950_ u_cpu.rf_ram_if.wdata1_r\[2\] net341 u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12793__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11321__A1 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11901_ _00423_ net90 u_cpu.rf_ram.memory\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12881_ _01378_ net507 u_cpu.rf_ram.memory\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11832_ _00354_ net12 u_cpu.rf_ram.memory\[68\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12023__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09817__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A1 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _00285_ net300 u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10714_ _04661_ _04777_ _04974_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11694_ _00216_ net402 u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10645_ _04068_ _05184_ _05187_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11388__A1 _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10576_ _05106_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12315_ _00816_ net485 u_cpu.rf_ram.memory\[35\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__A1 _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06091__I _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12246_ _00747_ net362 u_cpu.rf_ram.memory\[123\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08556__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12177_ _00691_ net425 u_cpu.rf_ram.memory\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10363__A2 _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11128_ u_cpu.rf_ram.memory\[69\]\[1\] _05502_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout198_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09505__A1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ _05399_ _05457_ _05459_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11312__A1 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09808__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout532_I net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12516__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ _03500_ _03526_ _03531_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07221_ _02749_ u_scanchain_local.module_data_in\[55\] _02788_ u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__A1 _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07152_ _02725_ _02727_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06103_ _01558_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09992__A1 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08795__A2 _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07083_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_dbus_dat\[22\] _02677_ _02679_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10516__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ _01537_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10452__S _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout104 net110 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout115 net117 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06558__A1 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11551__A1 _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout126 net130 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout137 net139 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout148 net150 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout159 net160 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07985_ u_cpu.rf_ram.memory\[40\]\[5\] _03338_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09724_ u_cpu.rf_ram.memory\[116\]\[5\] _04463_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06936_ _02573_ u_cpu.cpu.ctrl.i_iscomp _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10106__A2 _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09655_ u_cpu.rf_ram.memory\[112\]\[5\] _04418_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06867_ _01448_ _01449_ _01446_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_103_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _03751_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05818_ _01468_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08656__I _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09586_ _04337_ _04377_ _04380_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06730__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ _01730_ _02439_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08537_ _03550_ _03454_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12196__CLK net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10200__B _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06176__I _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _03581_ _03651_ _03660_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05916__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06333__I1 u_cpu.rf_ram.memory\[77\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ _02957_ _02959_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08399_ _03608_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10417__I0 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _05054_
+ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10361_ _02616_ _01441_ _04717_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06341__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10593__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12100_ _00614_ net260 u_cpu.rf_ram.memory\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10292_ u_cpu.cpu.immdec.imm19_12_20\[1\] _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12031_ _00545_ net420 u_cpu.rf_ram.memory\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09735__A1 u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06549__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11542__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10345__A2 _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12933_ _01429_ net379 u_cpu.rf_ram.memory\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06021__I0 u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08710__A2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12864_ _01361_ net500 u_cpu.rf_ram.memory\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11815_ _00337_ net18 u_cpu.rf_ram.memory\[75\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12795_ _01292_ net39 u_cpu.rf_ram.memory\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11746_ _00268_ net431 u_cpu.rf_ram.memory\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06086__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08474__A1 _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10281__A1 _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11677_ _00199_ net464 u_cpu.rf_ram.memory\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10628_ _04070_ _05172_ _05177_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07029__A2 _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06088__I0 u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__I2 u_cpu.rf_ram.memory\[78\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _05134_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10584__A2 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12229_ _00017_ net287 u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11533__A1 _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06689__C _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout482_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07201__A2 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ _03198_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06721_ _02188_ _02363_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _02491_ _02522_ _04283_ _04285_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06652_ u_cpu.rf_ram.memory\[4\]\[6\] u_cpu.rf_ram.memory\[5\]\[6\] u_cpu.rf_ram.memory\[6\]\[6\]
+ u_cpu.rf_ram.memory\[7\]\[6\] _01561_ _01897_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07380__I _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ u_cpu.rf_ram_if.rgnt _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06583_ _01919_ _02226_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08322_ _03511_ _03553_ _03562_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08465__A1 u_cpu.rf_ram.memory\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__I1 u_cpu.rf_ram.memory\[89\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10272__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ u_cpu.rf_ram.memory\[65\]\[4\] _03518_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10447__S _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10272__B2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ _02714_ _02773_ _02774_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08184_ u_cpu.rf_ram.memory\[68\]\[4\] _03473_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07135_ _02701_ u_scanchain_local.module_data_in\[40\] _02625_ u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06779__A1 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07066_ _02669_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06017_ _01650_ _01655_ _01658_ _01664_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_82_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10327__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09971__S _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ u_cpu.rf_ram.memory\[40\]\[1\] _03331_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06951__A1 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09707_ _04442_ _04448_ _04456_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06919_ _02521_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07899_ _02505_ _02864_ _02528_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _04079_ _04403_ _04411_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06703__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12831__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ _04339_ _04365_ _04370_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ _00122_ net415 u_cpu.rf_ram.memory\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07259__A2 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12580_ _01078_ net329 u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11531_ _03630_ _05754_ _05759_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11462_ _03050_ _03068_ _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__A1 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09956__A1 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10413_ u_cpu.cpu.alu.cmp_r _02869_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08759__A2 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11393_ _05628_ _05670_ _05676_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10344_ _04986_ _04997_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07431__A2 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10092__S _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ _04831_ _04665_ _04692_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10318__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11515__A1 _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12014_ _00528_ net43 u_cpu.rf_ram.memory\[141\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09184__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07195__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07195__B2 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout490 net492 net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_48_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12916_ _01413_ net176 u_cpu.rf_ram.memory\[100\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07414__B u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12847_ _01344_ net437 u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12778_ _01275_ net13 u_cpu.rf_ram.memory\[69\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout230_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__B2 u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08998__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11729_ _00251_ net219 u_cpu.rf_ram.memory\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout328_I net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10006__A1 _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09947__A1 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__S0 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06225__A3 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07422__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _03957_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11506__A1 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10309__A2 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05984__A2 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09175__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ _03848_ _03914_ _03917_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06608__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07186__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13029__D _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07822_ u_cpu.rf_ram.memory\[47\]\[0\] _03234_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08922__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06784__I1 u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ _03137_ _03185_ _03188_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06704_ u_cpu.rf_ram.memory\[80\]\[6\] u_cpu.rf_ram.memory\[81\]\[6\] u_cpu.rf_ram.memory\[82\]\[6\]
+ u_cpu.rf_ram.memory\[83\]\[6\] _01584_ _01965_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07489__A2 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _02927_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ _04258_ _04267_ _04274_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06635_ _01763_ _02278_ _01756_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06792__S0 _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09354_ u_cpu.rf_ram.memory\[36\]\[7\] _04216_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06566_ u_cpu.rf_ram.memory\[0\]\[5\] u_cpu.rf_ram.memory\[1\]\[5\] u_cpu.rf_ram.memory\[2\]\[5\]
+ u_cpu.rf_ram.memory\[3\]\[5\] _01786_ _01900_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08934__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08305_ _03551_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08989__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09285_ _04161_ _04181_ _04186_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06497_ u_cpu.rf_ram.memory\[52\]\[4\] u_cpu.rf_ram.memory\[53\]\[4\] u_cpu.rf_ram.memory\[54\]\[4\]
+ u_cpu.rf_ram.memory\[55\]\[4\] _01630_ _02040_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06544__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08236_ u_cpu.rf_ram.memory\[66\]\[6\] _03501_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12234__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07661__A2 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ _02940_ _03458_ _03465_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10548__A2 _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ _02621_ u_cpu.cpu.state.ibus_cyc _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _03420_ _03410_ _03421_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06472__I0 u_cpu.rf_ram.memory\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ u_arbiter.i_wb_cpu_rdt\[10\] u_arbiter.i_wb_cpu_dbus_dat\[7\] _02658_ _02660_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _04743_ _04721_ _04745_ _04703_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06924__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10962_ u_cpu.rf_ram.memory\[104\]\[6\] _05392_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06527__I1 u_cpu.rf_ram.memory\[81\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12701_ _01198_ net137 u_cpu.rf_ram.memory\[103\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10893_ u_cpu.rf_ram.memory\[101\]\[2\] _05355_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12632_ _01129_ net154 u_cpu.rf_ram.memory\[97\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12563_ _01061_ net309 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10787__A2 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11514_ u_cpu.rf_ram.memory\[100\]\[4\] _05746_ _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07652__A2 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12494_ _00995_ net240 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09929__A1 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11445_ u_cpu.rf_ram.memory\[24\]\[0\] _05707_ _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12727__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09675__I _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07404__A2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11376_ u_cpu.cpu.genblk3.csr.mstatus_mie _05638_ _05663_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10327_ _04972_ _04973_ _04681_ _04981_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11751__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12877__CLK net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10258_ _04862_ _04908_ _04754_ _04919_ _04745_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ _04620_ _04849_ _04857_ _04600_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10711__A2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout180_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12107__CLK net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06230__I3 u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout278_I net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09865__B1 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout445_I net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ _01583_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12257__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07891__A2 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06351_ _01497_ _01933_ _01997_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09093__A1 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10778__A2 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09070_ u_cpu.rf_ram.memory\[131\]\[2\] _04043_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06282_ _01595_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07643__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__A1 u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08021_ _03371_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__A2 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10250__I1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09972_ _04663_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07319__B _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08923_ u_cpu.rf_ram.memory\[137\]\[3\] _03950_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07159__A1 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08854_ _03631_ _03902_ _03907_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10163__B1 _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10702__A2 _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07805_ _02933_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _03863_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05997_ _01628_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07736_ u_cpu.rf_ram.memory\[51\]\[4\] _03174_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08659__A1 u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07667_ _03031_ _03119_ _03128_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ _04262_ _04249_ _04263_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06618_ u_cpu.rf_ram.memory\[84\]\[5\] u_cpu.rf_ram.memory\[85\]\[5\] u_cpu.rf_ram.memory\[86\]\[5\]
+ u_cpu.rf_ram.memory\[87\]\[5\] _01855_ _02083_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07598_ _03082_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_90_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__A1 _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06549_ _01758_ _02193_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09337_ _04216_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06517__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10769__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06184__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04173_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06288__I3 u_cpu.rf_ram.memory\[103\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ _03333_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09199_ _03082_ _03356_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11230_ _05220_ _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__A2 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11774__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07398__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11194__A2 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _05484_ _05515_ _05523_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05948__A2 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10941__A2 _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09139__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _04726_ _04793_ _04782_ _04624_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_27_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11092_ u_cpu.rf_ram.memory\[83\]\[4\] _05476_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10043_ _04721_ _04729_ _04704_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06212__I3 u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07570__A1 u_cpu.rf_ram.memory\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11994_ _00516_ net223 u_cpu.rf_ram.memory\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10945_ _05328_ _05377_ _05386_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06125__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07322__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__A2 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10876_ _04632_ _05331_ _05345_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12615_ _01112_ net159 u_cpu.rf_ram.memory\[93\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09075__A1 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06508__S0 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06308__B _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06094__I _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12546_ _01046_ net187 u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06428__A3 _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08822__A1 _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12477_ _00978_ net238 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07918__I _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11428_ _05623_ _05694_ _05697_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11359_ _02539_ _05643_ _05640_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05939__A2 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10932__A2 _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout395_I net397 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05920_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13029_ _00091_ net534 u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05851_ _01467_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10696__A1 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09550__A2 _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__A2 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08570_ _03673_ _03718_ _03725_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09838__B1 _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07521_ _02951_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_81_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11647__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _02984_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07864__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05901__I _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06403_ _01646_ _02048_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ u_cpu.rf_ram.memory\[82\]\[3\] _02922_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10519__I _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09066__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _02939_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06334_ _01735_ _01980_ _01738_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07616__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ _04003_ _04027_ _04033_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06265_ _01589_ _01911_ _01801_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08004_ _03357_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _01683_ _01843_ _01687_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11176__A2 _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__A2 _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _04602_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08906_ _03939_ _03928_ _03940_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09886_ _04584_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _03855_ _03889_ _03896_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06179__I _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09829__B1 _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _03742_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ u_cpu.rf_ram.memory\[44\]\[7\] _03154_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ u_cpu.rf_ram.memory\[140\]\[1\] _03808_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _04782_ _05253_ _04665_ _04791_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10661_ _04295_ _03132_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09057__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06128__B _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12400_ _00901_ net459 u_cpu.rf_ram.memory\[116\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _02577_ _02554_ u_cpu.cpu.ctrl.i_jump _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10611__A1 u_cpu.rf_ram.memory\[109\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12331_ _00832_ net454 u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10365__S _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__A2 _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12262_ _00763_ net360 u_cpu.rf_ram.memory\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06830__A3 u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11167__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11213_ _05555_ _05552_ _05556_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput6 net6 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_12193_ _00707_ net268 u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08032__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11144_ _05512_ _03013_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09780__A2 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11075_ _05195_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10678__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ _02708_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A2 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12915__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06089__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12966__D _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09296__A1 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11977_ _00499_ net58 u_cpu.rf_ram.memory\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _05375_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout143_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09048__A1 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10859_ _05336_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10602__A1 u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout310_I net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12529_ _01030_ net324 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout408_I net409 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08271__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ _01635_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08023__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__A2 _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout308 net312 net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout319 net320 net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06424__I3 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__A1 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__I _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09740_ u_cpu.rf_ram.memory\[33\]\[3\] _04475_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06952_ _02584_ _02586_ _02588_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

