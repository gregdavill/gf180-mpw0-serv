magic
tech gf180mcuC
magscale 1 5
timestamp 1670140657
<< obsm1 >>
rect 672 1538 69328 58438
<< metal2 >>
rect 2184 59800 2240 60000
rect 2744 59800 2800 60000
rect 3304 59800 3360 60000
rect 3864 59800 3920 60000
rect 4424 59800 4480 60000
rect 4984 59800 5040 60000
rect 5544 59800 5600 60000
rect 6104 59800 6160 60000
rect 6664 59800 6720 60000
rect 7224 59800 7280 60000
rect 7784 59800 7840 60000
rect 8344 59800 8400 60000
rect 8904 59800 8960 60000
rect 9464 59800 9520 60000
rect 10024 59800 10080 60000
rect 10584 59800 10640 60000
rect 11144 59800 11200 60000
rect 11704 59800 11760 60000
rect 12264 59800 12320 60000
rect 12824 59800 12880 60000
rect 13384 59800 13440 60000
rect 13944 59800 14000 60000
rect 14504 59800 14560 60000
rect 15064 59800 15120 60000
rect 15624 59800 15680 60000
rect 16184 59800 16240 60000
rect 16744 59800 16800 60000
rect 17304 59800 17360 60000
rect 17864 59800 17920 60000
rect 18424 59800 18480 60000
rect 18984 59800 19040 60000
rect 19544 59800 19600 60000
rect 20104 59800 20160 60000
rect 20664 59800 20720 60000
rect 21224 59800 21280 60000
rect 21784 59800 21840 60000
rect 22344 59800 22400 60000
rect 22904 59800 22960 60000
rect 23464 59800 23520 60000
rect 24024 59800 24080 60000
rect 24584 59800 24640 60000
rect 25144 59800 25200 60000
rect 25704 59800 25760 60000
rect 26264 59800 26320 60000
rect 26824 59800 26880 60000
rect 27384 59800 27440 60000
rect 27944 59800 28000 60000
rect 28504 59800 28560 60000
rect 29064 59800 29120 60000
rect 29624 59800 29680 60000
rect 30184 59800 30240 60000
rect 30744 59800 30800 60000
rect 31304 59800 31360 60000
rect 31864 59800 31920 60000
rect 32424 59800 32480 60000
rect 32984 59800 33040 60000
rect 33544 59800 33600 60000
rect 34104 59800 34160 60000
rect 34664 59800 34720 60000
rect 35224 59800 35280 60000
rect 35784 59800 35840 60000
rect 36344 59800 36400 60000
rect 36904 59800 36960 60000
rect 37464 59800 37520 60000
rect 38024 59800 38080 60000
rect 38584 59800 38640 60000
rect 39144 59800 39200 60000
rect 39704 59800 39760 60000
rect 40264 59800 40320 60000
rect 40824 59800 40880 60000
rect 41384 59800 41440 60000
rect 41944 59800 42000 60000
rect 42504 59800 42560 60000
rect 43064 59800 43120 60000
rect 43624 59800 43680 60000
rect 44184 59800 44240 60000
rect 44744 59800 44800 60000
rect 45304 59800 45360 60000
rect 45864 59800 45920 60000
rect 46424 59800 46480 60000
rect 46984 59800 47040 60000
rect 47544 59800 47600 60000
rect 48104 59800 48160 60000
rect 48664 59800 48720 60000
rect 49224 59800 49280 60000
rect 49784 59800 49840 60000
rect 50344 59800 50400 60000
rect 50904 59800 50960 60000
rect 51464 59800 51520 60000
rect 52024 59800 52080 60000
rect 52584 59800 52640 60000
rect 53144 59800 53200 60000
rect 53704 59800 53760 60000
rect 54264 59800 54320 60000
rect 54824 59800 54880 60000
rect 55384 59800 55440 60000
rect 55944 59800 56000 60000
rect 56504 59800 56560 60000
rect 57064 59800 57120 60000
rect 57624 59800 57680 60000
rect 58184 59800 58240 60000
rect 58744 59800 58800 60000
rect 59304 59800 59360 60000
rect 59864 59800 59920 60000
rect 60424 59800 60480 60000
rect 60984 59800 61040 60000
rect 61544 59800 61600 60000
rect 62104 59800 62160 60000
rect 62664 59800 62720 60000
rect 63224 59800 63280 60000
rect 63784 59800 63840 60000
rect 64344 59800 64400 60000
rect 64904 59800 64960 60000
rect 65464 59800 65520 60000
rect 66024 59800 66080 60000
rect 66584 59800 66640 60000
rect 67144 59800 67200 60000
rect 67704 59800 67760 60000
rect 1680 0 1736 200
rect 1904 0 1960 200
rect 2128 0 2184 200
rect 2352 0 2408 200
rect 2576 0 2632 200
rect 2800 0 2856 200
rect 3024 0 3080 200
rect 3248 0 3304 200
rect 3472 0 3528 200
rect 3696 0 3752 200
rect 3920 0 3976 200
rect 4144 0 4200 200
rect 4368 0 4424 200
rect 4592 0 4648 200
rect 4816 0 4872 200
rect 5040 0 5096 200
rect 5264 0 5320 200
rect 5488 0 5544 200
rect 5712 0 5768 200
rect 5936 0 5992 200
rect 6160 0 6216 200
rect 6384 0 6440 200
rect 6608 0 6664 200
rect 6832 0 6888 200
rect 7056 0 7112 200
rect 7280 0 7336 200
rect 7504 0 7560 200
rect 7728 0 7784 200
rect 7952 0 8008 200
rect 8176 0 8232 200
rect 8400 0 8456 200
rect 8624 0 8680 200
rect 8848 0 8904 200
rect 9072 0 9128 200
rect 9296 0 9352 200
rect 9520 0 9576 200
rect 9744 0 9800 200
rect 9968 0 10024 200
rect 10192 0 10248 200
rect 10416 0 10472 200
rect 10640 0 10696 200
rect 10864 0 10920 200
rect 11088 0 11144 200
rect 11312 0 11368 200
rect 11536 0 11592 200
rect 11760 0 11816 200
rect 11984 0 12040 200
rect 12208 0 12264 200
rect 12432 0 12488 200
rect 12656 0 12712 200
rect 12880 0 12936 200
rect 13104 0 13160 200
rect 13328 0 13384 200
rect 13552 0 13608 200
rect 13776 0 13832 200
rect 14000 0 14056 200
rect 14224 0 14280 200
rect 14448 0 14504 200
rect 14672 0 14728 200
rect 14896 0 14952 200
rect 15120 0 15176 200
rect 15344 0 15400 200
rect 15568 0 15624 200
rect 15792 0 15848 200
rect 16016 0 16072 200
rect 16240 0 16296 200
rect 16464 0 16520 200
rect 16688 0 16744 200
rect 16912 0 16968 200
rect 17136 0 17192 200
rect 17360 0 17416 200
rect 17584 0 17640 200
rect 17808 0 17864 200
rect 18032 0 18088 200
rect 18256 0 18312 200
rect 18480 0 18536 200
rect 18704 0 18760 200
rect 18928 0 18984 200
rect 19152 0 19208 200
rect 19376 0 19432 200
rect 19600 0 19656 200
rect 19824 0 19880 200
rect 20048 0 20104 200
rect 20272 0 20328 200
rect 20496 0 20552 200
rect 20720 0 20776 200
rect 20944 0 21000 200
rect 21168 0 21224 200
rect 21392 0 21448 200
rect 21616 0 21672 200
rect 21840 0 21896 200
rect 22064 0 22120 200
rect 22288 0 22344 200
rect 22512 0 22568 200
rect 22736 0 22792 200
rect 22960 0 23016 200
rect 23184 0 23240 200
rect 23408 0 23464 200
rect 23632 0 23688 200
rect 23856 0 23912 200
rect 24080 0 24136 200
rect 24304 0 24360 200
rect 24528 0 24584 200
rect 24752 0 24808 200
rect 24976 0 25032 200
rect 25200 0 25256 200
rect 25424 0 25480 200
rect 25648 0 25704 200
rect 25872 0 25928 200
rect 26096 0 26152 200
rect 26320 0 26376 200
rect 26544 0 26600 200
rect 26768 0 26824 200
rect 26992 0 27048 200
rect 27216 0 27272 200
rect 27440 0 27496 200
rect 27664 0 27720 200
rect 27888 0 27944 200
rect 28112 0 28168 200
rect 28336 0 28392 200
rect 28560 0 28616 200
rect 28784 0 28840 200
rect 29008 0 29064 200
rect 29232 0 29288 200
rect 29456 0 29512 200
rect 29680 0 29736 200
rect 29904 0 29960 200
rect 30128 0 30184 200
rect 30352 0 30408 200
rect 30576 0 30632 200
rect 30800 0 30856 200
rect 31024 0 31080 200
rect 31248 0 31304 200
rect 31472 0 31528 200
rect 31696 0 31752 200
rect 31920 0 31976 200
rect 32144 0 32200 200
rect 32368 0 32424 200
rect 32592 0 32648 200
rect 32816 0 32872 200
rect 33040 0 33096 200
rect 33264 0 33320 200
rect 33488 0 33544 200
rect 33712 0 33768 200
rect 33936 0 33992 200
rect 34160 0 34216 200
rect 34384 0 34440 200
rect 34608 0 34664 200
rect 34832 0 34888 200
rect 35056 0 35112 200
rect 35280 0 35336 200
rect 35504 0 35560 200
rect 35728 0 35784 200
rect 35952 0 36008 200
rect 36176 0 36232 200
rect 36400 0 36456 200
rect 36624 0 36680 200
rect 36848 0 36904 200
rect 37072 0 37128 200
rect 37296 0 37352 200
rect 37520 0 37576 200
rect 37744 0 37800 200
rect 37968 0 38024 200
rect 38192 0 38248 200
rect 38416 0 38472 200
rect 38640 0 38696 200
rect 38864 0 38920 200
rect 39088 0 39144 200
rect 39312 0 39368 200
rect 39536 0 39592 200
rect 39760 0 39816 200
rect 39984 0 40040 200
rect 40208 0 40264 200
rect 40432 0 40488 200
rect 40656 0 40712 200
rect 40880 0 40936 200
rect 41104 0 41160 200
rect 41328 0 41384 200
rect 41552 0 41608 200
rect 41776 0 41832 200
rect 42000 0 42056 200
rect 42224 0 42280 200
rect 42448 0 42504 200
rect 42672 0 42728 200
rect 42896 0 42952 200
rect 43120 0 43176 200
rect 43344 0 43400 200
rect 43568 0 43624 200
rect 43792 0 43848 200
rect 44016 0 44072 200
rect 44240 0 44296 200
rect 44464 0 44520 200
rect 44688 0 44744 200
rect 44912 0 44968 200
rect 45136 0 45192 200
rect 45360 0 45416 200
rect 45584 0 45640 200
rect 45808 0 45864 200
rect 46032 0 46088 200
rect 46256 0 46312 200
rect 46480 0 46536 200
rect 46704 0 46760 200
rect 46928 0 46984 200
rect 47152 0 47208 200
rect 47376 0 47432 200
rect 47600 0 47656 200
rect 47824 0 47880 200
rect 48048 0 48104 200
rect 48272 0 48328 200
rect 48496 0 48552 200
rect 48720 0 48776 200
rect 48944 0 49000 200
rect 49168 0 49224 200
rect 49392 0 49448 200
rect 49616 0 49672 200
rect 49840 0 49896 200
rect 50064 0 50120 200
rect 50288 0 50344 200
rect 50512 0 50568 200
rect 50736 0 50792 200
rect 50960 0 51016 200
rect 51184 0 51240 200
rect 51408 0 51464 200
rect 51632 0 51688 200
rect 51856 0 51912 200
rect 52080 0 52136 200
rect 52304 0 52360 200
rect 52528 0 52584 200
rect 52752 0 52808 200
rect 52976 0 53032 200
rect 53200 0 53256 200
rect 53424 0 53480 200
rect 53648 0 53704 200
rect 53872 0 53928 200
rect 54096 0 54152 200
rect 54320 0 54376 200
rect 54544 0 54600 200
rect 54768 0 54824 200
rect 54992 0 55048 200
rect 55216 0 55272 200
rect 55440 0 55496 200
rect 55664 0 55720 200
rect 55888 0 55944 200
rect 56112 0 56168 200
rect 56336 0 56392 200
rect 56560 0 56616 200
rect 56784 0 56840 200
rect 57008 0 57064 200
rect 57232 0 57288 200
rect 57456 0 57512 200
rect 57680 0 57736 200
rect 57904 0 57960 200
rect 58128 0 58184 200
rect 58352 0 58408 200
rect 58576 0 58632 200
rect 58800 0 58856 200
rect 59024 0 59080 200
rect 59248 0 59304 200
rect 59472 0 59528 200
rect 59696 0 59752 200
rect 59920 0 59976 200
rect 60144 0 60200 200
rect 60368 0 60424 200
rect 60592 0 60648 200
rect 60816 0 60872 200
rect 61040 0 61096 200
rect 61264 0 61320 200
rect 61488 0 61544 200
rect 61712 0 61768 200
rect 61936 0 61992 200
rect 62160 0 62216 200
rect 62384 0 62440 200
rect 62608 0 62664 200
rect 62832 0 62888 200
rect 63056 0 63112 200
rect 63280 0 63336 200
rect 63504 0 63560 200
rect 63728 0 63784 200
rect 63952 0 64008 200
rect 64176 0 64232 200
rect 64400 0 64456 200
rect 64624 0 64680 200
rect 64848 0 64904 200
rect 65072 0 65128 200
rect 65296 0 65352 200
rect 65520 0 65576 200
rect 65744 0 65800 200
rect 65968 0 66024 200
rect 66192 0 66248 200
rect 66416 0 66472 200
rect 66640 0 66696 200
rect 66864 0 66920 200
rect 67088 0 67144 200
rect 67312 0 67368 200
rect 67536 0 67592 200
rect 67760 0 67816 200
rect 67984 0 68040 200
rect 68208 0 68264 200
<< obsm2 >>
rect 2142 59770 2154 59800
rect 2270 59770 2714 59800
rect 2830 59770 3274 59800
rect 3390 59770 3834 59800
rect 3950 59770 4394 59800
rect 4510 59770 4954 59800
rect 5070 59770 5514 59800
rect 5630 59770 6074 59800
rect 6190 59770 6634 59800
rect 6750 59770 7194 59800
rect 7310 59770 7754 59800
rect 7870 59770 8314 59800
rect 8430 59770 8874 59800
rect 8990 59770 9434 59800
rect 9550 59770 9994 59800
rect 10110 59770 10554 59800
rect 10670 59770 11114 59800
rect 11230 59770 11674 59800
rect 11790 59770 12234 59800
rect 12350 59770 12794 59800
rect 12910 59770 13354 59800
rect 13470 59770 13914 59800
rect 14030 59770 14474 59800
rect 14590 59770 15034 59800
rect 15150 59770 15594 59800
rect 15710 59770 16154 59800
rect 16270 59770 16714 59800
rect 16830 59770 17274 59800
rect 17390 59770 17834 59800
rect 17950 59770 18394 59800
rect 18510 59770 18954 59800
rect 19070 59770 19514 59800
rect 19630 59770 20074 59800
rect 20190 59770 20634 59800
rect 20750 59770 21194 59800
rect 21310 59770 21754 59800
rect 21870 59770 22314 59800
rect 22430 59770 22874 59800
rect 22990 59770 23434 59800
rect 23550 59770 23994 59800
rect 24110 59770 24554 59800
rect 24670 59770 25114 59800
rect 25230 59770 25674 59800
rect 25790 59770 26234 59800
rect 26350 59770 26794 59800
rect 26910 59770 27354 59800
rect 27470 59770 27914 59800
rect 28030 59770 28474 59800
rect 28590 59770 29034 59800
rect 29150 59770 29594 59800
rect 29710 59770 30154 59800
rect 30270 59770 30714 59800
rect 30830 59770 31274 59800
rect 31390 59770 31834 59800
rect 31950 59770 32394 59800
rect 32510 59770 32954 59800
rect 33070 59770 33514 59800
rect 33630 59770 34074 59800
rect 34190 59770 34634 59800
rect 34750 59770 35194 59800
rect 35310 59770 35754 59800
rect 35870 59770 36314 59800
rect 36430 59770 36874 59800
rect 36990 59770 37434 59800
rect 37550 59770 37994 59800
rect 38110 59770 38554 59800
rect 38670 59770 39114 59800
rect 39230 59770 39674 59800
rect 39790 59770 40234 59800
rect 40350 59770 40794 59800
rect 40910 59770 41354 59800
rect 41470 59770 41914 59800
rect 42030 59770 42474 59800
rect 42590 59770 43034 59800
rect 43150 59770 43594 59800
rect 43710 59770 44154 59800
rect 44270 59770 44714 59800
rect 44830 59770 45274 59800
rect 45390 59770 45834 59800
rect 45950 59770 46394 59800
rect 46510 59770 46954 59800
rect 47070 59770 47514 59800
rect 47630 59770 48074 59800
rect 48190 59770 48634 59800
rect 48750 59770 49194 59800
rect 49310 59770 49754 59800
rect 49870 59770 50314 59800
rect 50430 59770 50874 59800
rect 50990 59770 51434 59800
rect 51550 59770 51994 59800
rect 52110 59770 52554 59800
rect 52670 59770 53114 59800
rect 53230 59770 53674 59800
rect 53790 59770 54234 59800
rect 54350 59770 54794 59800
rect 54910 59770 55354 59800
rect 55470 59770 55914 59800
rect 56030 59770 56474 59800
rect 56590 59770 57034 59800
rect 57150 59770 57594 59800
rect 57710 59770 58154 59800
rect 58270 59770 58714 59800
rect 58830 59770 59274 59800
rect 59390 59770 59834 59800
rect 59950 59770 60394 59800
rect 60510 59770 60954 59800
rect 61070 59770 61514 59800
rect 61630 59770 62074 59800
rect 62190 59770 62634 59800
rect 62750 59770 63194 59800
rect 63310 59770 63754 59800
rect 63870 59770 64314 59800
rect 64430 59770 64874 59800
rect 64990 59770 65434 59800
rect 65550 59770 65994 59800
rect 66110 59770 66554 59800
rect 66670 59770 67114 59800
rect 67230 59770 67674 59800
rect 67790 59770 69314 59800
rect 2142 230 69314 59770
rect 2214 200 2322 230
rect 2438 200 2546 230
rect 2662 200 2770 230
rect 2886 200 2994 230
rect 3110 200 3218 230
rect 3334 200 3442 230
rect 3558 200 3666 230
rect 3782 200 3890 230
rect 4006 200 4114 230
rect 4230 200 4338 230
rect 4454 200 4562 230
rect 4678 200 4786 230
rect 4902 200 5010 230
rect 5126 200 5234 230
rect 5350 200 5458 230
rect 5574 200 5682 230
rect 5798 200 5906 230
rect 6022 200 6130 230
rect 6246 200 6354 230
rect 6470 200 6578 230
rect 6694 200 6802 230
rect 6918 200 7026 230
rect 7142 200 7250 230
rect 7366 200 7474 230
rect 7590 200 7698 230
rect 7814 200 7922 230
rect 8038 200 8146 230
rect 8262 200 8370 230
rect 8486 200 8594 230
rect 8710 200 8818 230
rect 8934 200 9042 230
rect 9158 200 9266 230
rect 9382 200 9490 230
rect 9606 200 9714 230
rect 9830 200 9938 230
rect 10054 200 10162 230
rect 10278 200 10386 230
rect 10502 200 10610 230
rect 10726 200 10834 230
rect 10950 200 11058 230
rect 11174 200 11282 230
rect 11398 200 11506 230
rect 11622 200 11730 230
rect 11846 200 11954 230
rect 12070 200 12178 230
rect 12294 200 12402 230
rect 12518 200 12626 230
rect 12742 200 12850 230
rect 12966 200 13074 230
rect 13190 200 13298 230
rect 13414 200 13522 230
rect 13638 200 13746 230
rect 13862 200 13970 230
rect 14086 200 14194 230
rect 14310 200 14418 230
rect 14534 200 14642 230
rect 14758 200 14866 230
rect 14982 200 15090 230
rect 15206 200 15314 230
rect 15430 200 15538 230
rect 15654 200 15762 230
rect 15878 200 15986 230
rect 16102 200 16210 230
rect 16326 200 16434 230
rect 16550 200 16658 230
rect 16774 200 16882 230
rect 16998 200 17106 230
rect 17222 200 17330 230
rect 17446 200 17554 230
rect 17670 200 17778 230
rect 17894 200 18002 230
rect 18118 200 18226 230
rect 18342 200 18450 230
rect 18566 200 18674 230
rect 18790 200 18898 230
rect 19014 200 19122 230
rect 19238 200 19346 230
rect 19462 200 19570 230
rect 19686 200 19794 230
rect 19910 200 20018 230
rect 20134 200 20242 230
rect 20358 200 20466 230
rect 20582 200 20690 230
rect 20806 200 20914 230
rect 21030 200 21138 230
rect 21254 200 21362 230
rect 21478 200 21586 230
rect 21702 200 21810 230
rect 21926 200 22034 230
rect 22150 200 22258 230
rect 22374 200 22482 230
rect 22598 200 22706 230
rect 22822 200 22930 230
rect 23046 200 23154 230
rect 23270 200 23378 230
rect 23494 200 23602 230
rect 23718 200 23826 230
rect 23942 200 24050 230
rect 24166 200 24274 230
rect 24390 200 24498 230
rect 24614 200 24722 230
rect 24838 200 24946 230
rect 25062 200 25170 230
rect 25286 200 25394 230
rect 25510 200 25618 230
rect 25734 200 25842 230
rect 25958 200 26066 230
rect 26182 200 26290 230
rect 26406 200 26514 230
rect 26630 200 26738 230
rect 26854 200 26962 230
rect 27078 200 27186 230
rect 27302 200 27410 230
rect 27526 200 27634 230
rect 27750 200 27858 230
rect 27974 200 28082 230
rect 28198 200 28306 230
rect 28422 200 28530 230
rect 28646 200 28754 230
rect 28870 200 28978 230
rect 29094 200 29202 230
rect 29318 200 29426 230
rect 29542 200 29650 230
rect 29766 200 29874 230
rect 29990 200 30098 230
rect 30214 200 30322 230
rect 30438 200 30546 230
rect 30662 200 30770 230
rect 30886 200 30994 230
rect 31110 200 31218 230
rect 31334 200 31442 230
rect 31558 200 31666 230
rect 31782 200 31890 230
rect 32006 200 32114 230
rect 32230 200 32338 230
rect 32454 200 32562 230
rect 32678 200 32786 230
rect 32902 200 33010 230
rect 33126 200 33234 230
rect 33350 200 33458 230
rect 33574 200 33682 230
rect 33798 200 33906 230
rect 34022 200 34130 230
rect 34246 200 34354 230
rect 34470 200 34578 230
rect 34694 200 34802 230
rect 34918 200 35026 230
rect 35142 200 35250 230
rect 35366 200 35474 230
rect 35590 200 35698 230
rect 35814 200 35922 230
rect 36038 200 36146 230
rect 36262 200 36370 230
rect 36486 200 36594 230
rect 36710 200 36818 230
rect 36934 200 37042 230
rect 37158 200 37266 230
rect 37382 200 37490 230
rect 37606 200 37714 230
rect 37830 200 37938 230
rect 38054 200 38162 230
rect 38278 200 38386 230
rect 38502 200 38610 230
rect 38726 200 38834 230
rect 38950 200 39058 230
rect 39174 200 39282 230
rect 39398 200 39506 230
rect 39622 200 39730 230
rect 39846 200 39954 230
rect 40070 200 40178 230
rect 40294 200 40402 230
rect 40518 200 40626 230
rect 40742 200 40850 230
rect 40966 200 41074 230
rect 41190 200 41298 230
rect 41414 200 41522 230
rect 41638 200 41746 230
rect 41862 200 41970 230
rect 42086 200 42194 230
rect 42310 200 42418 230
rect 42534 200 42642 230
rect 42758 200 42866 230
rect 42982 200 43090 230
rect 43206 200 43314 230
rect 43430 200 43538 230
rect 43654 200 43762 230
rect 43878 200 43986 230
rect 44102 200 44210 230
rect 44326 200 44434 230
rect 44550 200 44658 230
rect 44774 200 44882 230
rect 44998 200 45106 230
rect 45222 200 45330 230
rect 45446 200 45554 230
rect 45670 200 45778 230
rect 45894 200 46002 230
rect 46118 200 46226 230
rect 46342 200 46450 230
rect 46566 200 46674 230
rect 46790 200 46898 230
rect 47014 200 47122 230
rect 47238 200 47346 230
rect 47462 200 47570 230
rect 47686 200 47794 230
rect 47910 200 48018 230
rect 48134 200 48242 230
rect 48358 200 48466 230
rect 48582 200 48690 230
rect 48806 200 48914 230
rect 49030 200 49138 230
rect 49254 200 49362 230
rect 49478 200 49586 230
rect 49702 200 49810 230
rect 49926 200 50034 230
rect 50150 200 50258 230
rect 50374 200 50482 230
rect 50598 200 50706 230
rect 50822 200 50930 230
rect 51046 200 51154 230
rect 51270 200 51378 230
rect 51494 200 51602 230
rect 51718 200 51826 230
rect 51942 200 52050 230
rect 52166 200 52274 230
rect 52390 200 52498 230
rect 52614 200 52722 230
rect 52838 200 52946 230
rect 53062 200 53170 230
rect 53286 200 53394 230
rect 53510 200 53618 230
rect 53734 200 53842 230
rect 53958 200 54066 230
rect 54182 200 54290 230
rect 54406 200 54514 230
rect 54630 200 54738 230
rect 54854 200 54962 230
rect 55078 200 55186 230
rect 55302 200 55410 230
rect 55526 200 55634 230
rect 55750 200 55858 230
rect 55974 200 56082 230
rect 56198 200 56306 230
rect 56422 200 56530 230
rect 56646 200 56754 230
rect 56870 200 56978 230
rect 57094 200 57202 230
rect 57318 200 57426 230
rect 57542 200 57650 230
rect 57766 200 57874 230
rect 57990 200 58098 230
rect 58214 200 58322 230
rect 58438 200 58546 230
rect 58662 200 58770 230
rect 58886 200 58994 230
rect 59110 200 59218 230
rect 59334 200 59442 230
rect 59558 200 59666 230
rect 59782 200 59890 230
rect 60006 200 60114 230
rect 60230 200 60338 230
rect 60454 200 60562 230
rect 60678 200 60786 230
rect 60902 200 61010 230
rect 61126 200 61234 230
rect 61350 200 61458 230
rect 61574 200 61682 230
rect 61798 200 61906 230
rect 62022 200 62130 230
rect 62246 200 62354 230
rect 62470 200 62578 230
rect 62694 200 62802 230
rect 62918 200 63026 230
rect 63142 200 63250 230
rect 63366 200 63474 230
rect 63590 200 63698 230
rect 63814 200 63922 230
rect 64038 200 64146 230
rect 64262 200 64370 230
rect 64486 200 64594 230
rect 64710 200 64818 230
rect 64934 200 65042 230
rect 65158 200 65266 230
rect 65382 200 65490 230
rect 65606 200 65714 230
rect 65830 200 65938 230
rect 66054 200 66162 230
rect 66278 200 66386 230
rect 66502 200 66610 230
rect 66726 200 66834 230
rect 66950 200 67058 230
rect 67174 200 67282 230
rect 67398 200 67506 230
rect 67622 200 67730 230
rect 67846 200 67954 230
rect 68070 200 68178 230
rect 68294 200 69314 230
<< obsm3 >>
rect 2233 1554 69319 58422
<< metal4 >>
rect 2224 1538 2384 58438
rect 3724 1538 3884 58438
rect 5224 1538 5384 58438
rect 6724 1538 6884 58438
rect 8224 1538 8384 58438
rect 9724 1538 9884 58438
rect 11224 1538 11384 58438
rect 12724 1538 12884 58438
rect 14224 1538 14384 58438
rect 15724 1538 15884 58438
rect 17224 1538 17384 58438
rect 18724 1538 18884 58438
rect 20224 1538 20384 58438
rect 21724 1538 21884 58438
rect 23224 1538 23384 58438
rect 24724 1538 24884 58438
rect 26224 1538 26384 58438
rect 27724 1538 27884 58438
rect 29224 1538 29384 58438
rect 30724 1538 30884 58438
rect 32224 1538 32384 58438
rect 33724 1538 33884 58438
rect 35224 1538 35384 58438
rect 36724 1538 36884 58438
rect 38224 1538 38384 58438
rect 39724 1538 39884 58438
rect 41224 1538 41384 58438
rect 42724 1538 42884 58438
rect 44224 1538 44384 58438
rect 45724 1538 45884 58438
rect 47224 1538 47384 58438
rect 48724 1538 48884 58438
rect 50224 1538 50384 58438
rect 51724 1538 51884 58438
rect 53224 1538 53384 58438
rect 54724 1538 54884 58438
rect 56224 1538 56384 58438
rect 57724 1538 57884 58438
rect 59224 1538 59384 58438
rect 60724 1538 60884 58438
rect 62224 1538 62384 58438
rect 63724 1538 63884 58438
rect 65224 1538 65384 58438
rect 66724 1538 66884 58438
rect 68224 1538 68384 58438
<< obsm4 >>
rect 34566 6337 35194 40647
rect 35414 6337 36694 40647
rect 36914 6337 38194 40647
rect 38414 6337 39694 40647
rect 39914 6337 41194 40647
rect 41414 6337 42694 40647
rect 42914 6337 44194 40647
rect 44414 6337 45694 40647
rect 45914 6337 47194 40647
rect 47414 6337 48694 40647
rect 48914 6337 50194 40647
rect 50414 6337 51694 40647
rect 51914 6337 53194 40647
rect 53414 6337 54694 40647
rect 54914 6337 56194 40647
rect 56414 6337 57694 40647
rect 57914 6337 59194 40647
rect 59414 6337 60694 40647
rect 60914 6337 62194 40647
rect 62414 6337 63694 40647
rect 63914 6337 65194 40647
rect 65414 6337 66694 40647
rect 66914 6337 68194 40647
rect 68414 6337 68978 40647
<< labels >>
rlabel metal2 s 2184 59800 2240 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 18984 59800 19040 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 20664 59800 20720 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 22344 59800 22400 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 24024 59800 24080 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 25704 59800 25760 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 27384 59800 27440 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 29064 59800 29120 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 30744 59800 30800 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 32424 59800 32480 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 34104 59800 34160 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3864 59800 3920 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 35784 59800 35840 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 37464 59800 37520 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 39144 59800 39200 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 40824 59800 40880 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 42504 59800 42560 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 44184 59800 44240 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 45864 59800 45920 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 47544 59800 47600 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 49224 59800 49280 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 50904 59800 50960 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5544 59800 5600 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 52584 59800 52640 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 54264 59800 54320 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 55944 59800 56000 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 57624 59800 57680 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 59304 59800 59360 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 60984 59800 61040 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 62664 59800 62720 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 64344 59800 64400 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7224 59800 7280 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 8904 59800 8960 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 10584 59800 10640 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 12264 59800 12320 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 13944 59800 14000 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 15624 59800 15680 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 17304 59800 17360 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2744 59800 2800 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 19544 59800 19600 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 21224 59800 21280 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 22904 59800 22960 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 24584 59800 24640 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 26264 59800 26320 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 27944 59800 28000 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 29624 59800 29680 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 31304 59800 31360 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 32984 59800 33040 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 34664 59800 34720 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4424 59800 4480 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 36344 59800 36400 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 38024 59800 38080 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 39704 59800 39760 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 41384 59800 41440 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 43064 59800 43120 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 44744 59800 44800 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 46424 59800 46480 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 48104 59800 48160 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 49784 59800 49840 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 51464 59800 51520 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6104 59800 6160 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 53144 59800 53200 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 54824 59800 54880 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 56504 59800 56560 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 58184 59800 58240 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 59864 59800 59920 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 61544 59800 61600 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 63224 59800 63280 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 64904 59800 64960 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 7784 59800 7840 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 9464 59800 9520 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 11144 59800 11200 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 12824 59800 12880 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 14504 59800 14560 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 16184 59800 16240 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 17864 59800 17920 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3304 59800 3360 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 20104 59800 20160 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 21784 59800 21840 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 23464 59800 23520 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 25144 59800 25200 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 26824 59800 26880 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 28504 59800 28560 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 30184 59800 30240 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 31864 59800 31920 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 33544 59800 33600 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 35224 59800 35280 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4984 59800 5040 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 36904 59800 36960 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 38584 59800 38640 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 40264 59800 40320 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 41944 59800 42000 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 43624 59800 43680 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 45304 59800 45360 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 46984 59800 47040 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 48664 59800 48720 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 50344 59800 50400 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 52024 59800 52080 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6664 59800 6720 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 53704 59800 53760 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 55384 59800 55440 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 57064 59800 57120 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 58744 59800 58800 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 60424 59800 60480 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 62104 59800 62160 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 63784 59800 63840 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 65464 59800 65520 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 8344 59800 8400 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 10024 59800 10080 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 11704 59800 11760 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 13384 59800 13440 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 15064 59800 15120 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 16744 59800 16800 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 18424 59800 18480 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 25424 0 25480 200 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 32144 0 32200 200 6 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 32816 0 32872 200 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 33488 0 33544 200 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 34160 0 34216 200 6 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 34832 0 34888 200 6 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 35504 0 35560 200 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 36176 0 36232 200 6 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 36848 0 36904 200 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 37520 0 37576 200 6 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 38192 0 38248 200 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 26096 0 26152 200 6 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 38864 0 38920 200 6 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 39536 0 39592 200 6 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 40208 0 40264 200 6 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 40880 0 40936 200 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 41552 0 41608 200 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 42224 0 42280 200 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 42896 0 42952 200 6 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 43568 0 43624 200 6 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 44240 0 44296 200 6 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 44912 0 44968 200 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 26768 0 26824 200 6 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 45584 0 45640 200 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 46256 0 46312 200 6 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 46928 0 46984 200 6 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 47600 0 47656 200 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 48272 0 48328 200 6 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 48944 0 49000 200 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 49616 0 49672 200 6 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 50288 0 50344 200 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 50960 0 51016 200 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 51632 0 51688 200 6 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 27440 0 27496 200 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 52304 0 52360 200 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 52976 0 53032 200 6 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 53648 0 53704 200 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 54320 0 54376 200 6 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 54992 0 55048 200 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 55664 0 55720 200 6 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 56336 0 56392 200 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 57008 0 57064 200 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 57680 0 57736 200 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 58352 0 58408 200 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 28112 0 28168 200 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 59024 0 59080 200 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 59696 0 59752 200 6 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 60368 0 60424 200 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 61040 0 61096 200 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 61712 0 61768 200 6 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 62384 0 62440 200 6 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 63056 0 63112 200 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 63728 0 63784 200 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 64400 0 64456 200 6 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 65072 0 65128 200 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 28784 0 28840 200 6 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 65744 0 65800 200 6 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 66416 0 66472 200 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 67088 0 67144 200 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 67760 0 67816 200 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 29456 0 29512 200 6 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 30128 0 30184 200 6 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 30800 0 30856 200 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 31472 0 31528 200 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 25648 0 25704 200 6 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 32368 0 32424 200 6 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 33040 0 33096 200 6 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 33712 0 33768 200 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 34384 0 34440 200 6 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 35056 0 35112 200 6 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 35728 0 35784 200 6 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 36400 0 36456 200 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 37072 0 37128 200 6 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 37744 0 37800 200 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 38416 0 38472 200 6 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 26320 0 26376 200 6 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 39088 0 39144 200 6 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 39760 0 39816 200 6 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 40432 0 40488 200 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 41104 0 41160 200 6 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 41776 0 41832 200 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 42448 0 42504 200 6 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 43120 0 43176 200 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 43792 0 43848 200 6 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 44464 0 44520 200 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 45136 0 45192 200 6 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 26992 0 27048 200 6 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 45808 0 45864 200 6 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 46480 0 46536 200 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 47152 0 47208 200 6 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 47824 0 47880 200 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 48496 0 48552 200 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 49168 0 49224 200 6 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 49840 0 49896 200 6 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 50512 0 50568 200 6 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 51184 0 51240 200 6 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 51856 0 51912 200 6 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 27664 0 27720 200 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 52528 0 52584 200 6 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 53200 0 53256 200 6 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 53872 0 53928 200 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 54544 0 54600 200 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 55216 0 55272 200 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 55888 0 55944 200 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 56560 0 56616 200 6 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 57232 0 57288 200 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 57904 0 57960 200 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 58576 0 58632 200 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 28336 0 28392 200 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 59248 0 59304 200 6 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 59920 0 59976 200 6 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 60592 0 60648 200 6 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 61264 0 61320 200 6 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 61936 0 61992 200 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 62608 0 62664 200 6 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 63280 0 63336 200 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 63952 0 64008 200 6 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 64624 0 64680 200 6 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 65296 0 65352 200 6 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 29008 0 29064 200 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 65968 0 66024 200 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 66640 0 66696 200 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 67312 0 67368 200 6 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 67984 0 68040 200 6 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 29680 0 29736 200 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 30352 0 30408 200 6 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 31024 0 31080 200 6 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 31696 0 31752 200 6 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 25872 0 25928 200 6 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 32592 0 32648 200 6 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 33264 0 33320 200 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 33936 0 33992 200 6 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 34608 0 34664 200 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 35280 0 35336 200 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 35952 0 36008 200 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 36624 0 36680 200 6 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 37296 0 37352 200 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 37968 0 38024 200 6 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 38640 0 38696 200 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 26544 0 26600 200 6 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 39312 0 39368 200 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 39984 0 40040 200 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 40656 0 40712 200 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 41328 0 41384 200 6 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 42000 0 42056 200 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 42672 0 42728 200 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 43344 0 43400 200 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 44016 0 44072 200 6 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 44688 0 44744 200 6 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 45360 0 45416 200 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 27216 0 27272 200 6 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 46032 0 46088 200 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 46704 0 46760 200 6 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 47376 0 47432 200 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 48048 0 48104 200 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 48720 0 48776 200 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 49392 0 49448 200 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 50064 0 50120 200 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 50736 0 50792 200 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 51408 0 51464 200 6 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 52080 0 52136 200 6 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 27888 0 27944 200 6 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 52752 0 52808 200 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 53424 0 53480 200 6 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 54096 0 54152 200 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 54768 0 54824 200 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 55440 0 55496 200 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 56112 0 56168 200 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 56784 0 56840 200 6 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 57456 0 57512 200 6 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 58128 0 58184 200 6 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 58800 0 58856 200 6 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 28560 0 28616 200 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 59472 0 59528 200 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 60144 0 60200 200 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 60816 0 60872 200 6 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 61488 0 61544 200 6 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 62160 0 62216 200 6 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 62832 0 62888 200 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 63504 0 63560 200 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 64176 0 64232 200 6 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 64848 0 64904 200 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 65520 0 65576 200 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 29232 0 29288 200 6 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 66192 0 66248 200 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 66864 0 66920 200 6 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 67536 0 67592 200 6 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 68208 0 68264 200 6 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 29904 0 29960 200 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 30576 0 30632 200 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 31248 0 31304 200 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 31920 0 31976 200 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 66024 59800 66080 60000 6 user_clock2
port 307 nsew signal input
rlabel metal2 s 66584 59800 66640 60000 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 67144 59800 67200 60000 6 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 67704 59800 67760 60000 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 5224 1538 5384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 8224 1538 8384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 11224 1538 11384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 14224 1538 14384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17224 1538 17384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 20224 1538 20384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 23224 1538 23384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 26224 1538 26384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 29224 1538 29384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32224 1538 32384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 35224 1538 35384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 38224 1538 38384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 41224 1538 41384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 44224 1538 44384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 47224 1538 47384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 50224 1538 50384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 53224 1538 53384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 56224 1538 56384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 59224 1538 59384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 62224 1538 62384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 65224 1538 65384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 68224 1538 68384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 3724 1538 3884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 6724 1538 6884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 9724 1538 9884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 12724 1538 12884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 15724 1538 15884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 18724 1538 18884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 21724 1538 21884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 24724 1538 24884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 27724 1538 27884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 30724 1538 30884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 33724 1538 33884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 36724 1538 36884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 39724 1538 39884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 42724 1538 42884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 45724 1538 45884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 48724 1538 48884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 51724 1538 51884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 54724 1538 54884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 57724 1538 57884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 60724 1538 60884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 63724 1538 63884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 66724 1538 66884 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 1680 0 1736 200 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 1904 0 1960 200 6 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 2128 0 2184 200 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 3024 0 3080 200 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 10640 0 10696 200 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 11312 0 11368 200 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 11984 0 12040 200 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 12656 0 12712 200 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 13328 0 13384 200 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 14000 0 14056 200 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 14672 0 14728 200 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 15344 0 15400 200 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 16016 0 16072 200 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 16688 0 16744 200 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 3920 0 3976 200 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 17360 0 17416 200 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 18032 0 18088 200 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 18704 0 18760 200 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 19376 0 19432 200 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 20048 0 20104 200 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 20720 0 20776 200 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 21392 0 21448 200 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 22064 0 22120 200 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 22736 0 22792 200 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 23408 0 23464 200 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 4816 0 4872 200 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 24080 0 24136 200 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 24752 0 24808 200 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 5712 0 5768 200 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 6608 0 6664 200 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 7280 0 7336 200 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 7952 0 8008 200 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 8624 0 8680 200 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 9296 0 9352 200 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 9968 0 10024 200 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 2352 0 2408 200 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 3248 0 3304 200 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 10864 0 10920 200 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 11536 0 11592 200 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 12208 0 12264 200 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 12880 0 12936 200 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 13552 0 13608 200 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 14224 0 14280 200 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 14896 0 14952 200 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 15568 0 15624 200 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 16240 0 16296 200 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 16912 0 16968 200 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 4144 0 4200 200 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 17584 0 17640 200 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 18256 0 18312 200 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 18928 0 18984 200 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 19600 0 19656 200 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 20272 0 20328 200 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 20944 0 21000 200 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 21616 0 21672 200 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 22288 0 22344 200 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 22960 0 23016 200 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 23632 0 23688 200 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 5040 0 5096 200 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 24304 0 24360 200 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 24976 0 25032 200 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 5936 0 5992 200 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 6832 0 6888 200 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 7504 0 7560 200 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 8176 0 8232 200 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 8848 0 8904 200 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 9520 0 9576 200 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 10192 0 10248 200 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 3472 0 3528 200 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 11088 0 11144 200 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 11760 0 11816 200 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 12432 0 12488 200 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 13104 0 13160 200 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 13776 0 13832 200 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 14448 0 14504 200 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 15120 0 15176 200 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 15792 0 15848 200 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 16464 0 16520 200 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 17136 0 17192 200 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 4368 0 4424 200 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 17808 0 17864 200 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 18480 0 18536 200 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 19152 0 19208 200 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 19824 0 19880 200 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 20496 0 20552 200 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 21168 0 21224 200 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 21840 0 21896 200 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 22512 0 22568 200 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 23184 0 23240 200 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 23856 0 23912 200 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 5264 0 5320 200 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 24528 0 24584 200 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 25200 0 25256 200 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 6160 0 6216 200 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 7056 0 7112 200 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 7728 0 7784 200 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 8400 0 8456 200 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 9072 0 9128 200 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 9744 0 9800 200 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 10416 0 10472 200 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 3696 0 3752 200 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 4592 0 4648 200 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 5488 0 5544 200 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 6384 0 6440 200 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 2576 0 2632 200 6 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 2800 0 2856 200 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8762770
string GDS_FILE /home/runner/work/gf180-mpw0-serv/gf180-mpw0-serv/openlane/tiny_user_project/runs/22_12_04_07_54/results/signoff/tiny_user_project.magic.gds
string GDS_START 2661780
<< end >>

