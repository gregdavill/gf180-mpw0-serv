// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire net9;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net10;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net11;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net47;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net48;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net49;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net82;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net83;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net84;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net85;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net86;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net87;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire \mod.cpu.alu.add_cy_r ;
 wire \mod.cpu.alu.cmp_r ;
 wire \mod.cpu.alu.i_rs1 ;
 wire \mod.cpu.bne_or_bge ;
 wire \mod.cpu.branch_op ;
 wire \mod.cpu.bufreg.c_r ;
 wire \mod.cpu.bufreg.data[10] ;
 wire \mod.cpu.bufreg.data[11] ;
 wire \mod.cpu.bufreg.data[12] ;
 wire \mod.cpu.bufreg.data[13] ;
 wire \mod.cpu.bufreg.data[14] ;
 wire \mod.cpu.bufreg.data[15] ;
 wire \mod.cpu.bufreg.data[16] ;
 wire \mod.cpu.bufreg.data[17] ;
 wire \mod.cpu.bufreg.data[18] ;
 wire \mod.cpu.bufreg.data[19] ;
 wire \mod.cpu.bufreg.data[20] ;
 wire \mod.cpu.bufreg.data[21] ;
 wire \mod.cpu.bufreg.data[22] ;
 wire \mod.cpu.bufreg.data[23] ;
 wire \mod.cpu.bufreg.data[24] ;
 wire \mod.cpu.bufreg.data[25] ;
 wire \mod.cpu.bufreg.data[26] ;
 wire \mod.cpu.bufreg.data[27] ;
 wire \mod.cpu.bufreg.data[28] ;
 wire \mod.cpu.bufreg.data[29] ;
 wire \mod.cpu.bufreg.data[2] ;
 wire \mod.cpu.bufreg.data[30] ;
 wire \mod.cpu.bufreg.data[31] ;
 wire \mod.cpu.bufreg.data[3] ;
 wire \mod.cpu.bufreg.data[4] ;
 wire \mod.cpu.bufreg.data[5] ;
 wire \mod.cpu.bufreg.data[6] ;
 wire \mod.cpu.bufreg.data[7] ;
 wire \mod.cpu.bufreg.data[8] ;
 wire \mod.cpu.bufreg.data[9] ;
 wire \mod.cpu.bufreg.i_sh_signed ;
 wire \mod.cpu.bufreg.lsb[0] ;
 wire \mod.cpu.bufreg.lsb[1] ;
 wire \mod.cpu.bufreg2.dat[0] ;
 wire \mod.cpu.bufreg2.dat[10] ;
 wire \mod.cpu.bufreg2.dat[11] ;
 wire \mod.cpu.bufreg2.dat[12] ;
 wire \mod.cpu.bufreg2.dat[13] ;
 wire \mod.cpu.bufreg2.dat[14] ;
 wire \mod.cpu.bufreg2.dat[15] ;
 wire \mod.cpu.bufreg2.dat[16] ;
 wire \mod.cpu.bufreg2.dat[17] ;
 wire \mod.cpu.bufreg2.dat[18] ;
 wire \mod.cpu.bufreg2.dat[19] ;
 wire \mod.cpu.bufreg2.dat[1] ;
 wire \mod.cpu.bufreg2.dat[20] ;
 wire \mod.cpu.bufreg2.dat[21] ;
 wire \mod.cpu.bufreg2.dat[22] ;
 wire \mod.cpu.bufreg2.dat[23] ;
 wire \mod.cpu.bufreg2.dat[24] ;
 wire \mod.cpu.bufreg2.dat[25] ;
 wire \mod.cpu.bufreg2.dat[26] ;
 wire \mod.cpu.bufreg2.dat[27] ;
 wire \mod.cpu.bufreg2.dat[28] ;
 wire \mod.cpu.bufreg2.dat[29] ;
 wire \mod.cpu.bufreg2.dat[2] ;
 wire \mod.cpu.bufreg2.dat[30] ;
 wire \mod.cpu.bufreg2.dat[31] ;
 wire \mod.cpu.bufreg2.dat[3] ;
 wire \mod.cpu.bufreg2.dat[4] ;
 wire \mod.cpu.bufreg2.dat[5] ;
 wire \mod.cpu.bufreg2.dat[6] ;
 wire \mod.cpu.bufreg2.dat[7] ;
 wire \mod.cpu.bufreg2.dat[8] ;
 wire \mod.cpu.bufreg2.dat[9] ;
 wire \mod.cpu.bufreg2.i_cnt_done ;
 wire \mod.cpu.bufreg2.i_dat[0] ;
 wire \mod.cpu.bufreg2.i_dat[10] ;
 wire \mod.cpu.bufreg2.i_dat[11] ;
 wire \mod.cpu.bufreg2.i_dat[12] ;
 wire \mod.cpu.bufreg2.i_dat[13] ;
 wire \mod.cpu.bufreg2.i_dat[14] ;
 wire \mod.cpu.bufreg2.i_dat[15] ;
 wire \mod.cpu.bufreg2.i_dat[16] ;
 wire \mod.cpu.bufreg2.i_dat[17] ;
 wire \mod.cpu.bufreg2.i_dat[18] ;
 wire \mod.cpu.bufreg2.i_dat[19] ;
 wire \mod.cpu.bufreg2.i_dat[1] ;
 wire \mod.cpu.bufreg2.i_dat[20] ;
 wire \mod.cpu.bufreg2.i_dat[21] ;
 wire \mod.cpu.bufreg2.i_dat[22] ;
 wire \mod.cpu.bufreg2.i_dat[23] ;
 wire \mod.cpu.bufreg2.i_dat[24] ;
 wire \mod.cpu.bufreg2.i_dat[25] ;
 wire \mod.cpu.bufreg2.i_dat[26] ;
 wire \mod.cpu.bufreg2.i_dat[27] ;
 wire \mod.cpu.bufreg2.i_dat[28] ;
 wire \mod.cpu.bufreg2.i_dat[29] ;
 wire \mod.cpu.bufreg2.i_dat[2] ;
 wire \mod.cpu.bufreg2.i_dat[30] ;
 wire \mod.cpu.bufreg2.i_dat[31] ;
 wire \mod.cpu.bufreg2.i_dat[3] ;
 wire \mod.cpu.bufreg2.i_dat[4] ;
 wire \mod.cpu.bufreg2.i_dat[5] ;
 wire \mod.cpu.bufreg2.i_dat[6] ;
 wire \mod.cpu.bufreg2.i_dat[7] ;
 wire \mod.cpu.bufreg2.i_dat[8] ;
 wire \mod.cpu.bufreg2.i_dat[9] ;
 wire \mod.cpu.bufreg2.i_op_b_sel ;
 wire \mod.cpu.bufreg2.i_rs2 ;
 wire \mod.cpu.csr_d_sel ;
 wire \mod.cpu.csr_imm ;
 wire \mod.cpu.ctrl.i_jump ;
 wire \mod.cpu.ctrl.o_ibus_adr[0] ;
 wire \mod.cpu.ctrl.o_ibus_adr[10] ;
 wire \mod.cpu.ctrl.o_ibus_adr[11] ;
 wire \mod.cpu.ctrl.o_ibus_adr[12] ;
 wire \mod.cpu.ctrl.o_ibus_adr[13] ;
 wire \mod.cpu.ctrl.o_ibus_adr[14] ;
 wire \mod.cpu.ctrl.o_ibus_adr[15] ;
 wire \mod.cpu.ctrl.o_ibus_adr[16] ;
 wire \mod.cpu.ctrl.o_ibus_adr[17] ;
 wire \mod.cpu.ctrl.o_ibus_adr[18] ;
 wire \mod.cpu.ctrl.o_ibus_adr[19] ;
 wire \mod.cpu.ctrl.o_ibus_adr[1] ;
 wire \mod.cpu.ctrl.o_ibus_adr[20] ;
 wire \mod.cpu.ctrl.o_ibus_adr[21] ;
 wire \mod.cpu.ctrl.o_ibus_adr[22] ;
 wire \mod.cpu.ctrl.o_ibus_adr[23] ;
 wire \mod.cpu.ctrl.o_ibus_adr[24] ;
 wire \mod.cpu.ctrl.o_ibus_adr[25] ;
 wire \mod.cpu.ctrl.o_ibus_adr[26] ;
 wire \mod.cpu.ctrl.o_ibus_adr[27] ;
 wire \mod.cpu.ctrl.o_ibus_adr[28] ;
 wire \mod.cpu.ctrl.o_ibus_adr[29] ;
 wire \mod.cpu.ctrl.o_ibus_adr[2] ;
 wire \mod.cpu.ctrl.o_ibus_adr[30] ;
 wire \mod.cpu.ctrl.o_ibus_adr[31] ;
 wire \mod.cpu.ctrl.o_ibus_adr[3] ;
 wire \mod.cpu.ctrl.o_ibus_adr[4] ;
 wire \mod.cpu.ctrl.o_ibus_adr[5] ;
 wire \mod.cpu.ctrl.o_ibus_adr[6] ;
 wire \mod.cpu.ctrl.o_ibus_adr[7] ;
 wire \mod.cpu.ctrl.o_ibus_adr[8] ;
 wire \mod.cpu.ctrl.o_ibus_adr[9] ;
 wire \mod.cpu.ctrl.pc_plus_4_cy_r ;
 wire \mod.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \mod.cpu.decode.co_ebreak ;
 wire \mod.cpu.decode.co_mem_word ;
 wire \mod.cpu.decode.opcode[0] ;
 wire \mod.cpu.decode.opcode[1] ;
 wire \mod.cpu.decode.opcode[2] ;
 wire \mod.cpu.i_rf_ready ;
 wire \mod.cpu.i_timer_irq ;
 wire \mod.cpu.immdec.imm11_7[0] ;
 wire \mod.cpu.immdec.imm11_7[1] ;
 wire \mod.cpu.immdec.imm11_7[2] ;
 wire \mod.cpu.immdec.imm11_7[3] ;
 wire \mod.cpu.immdec.imm11_7[4] ;
 wire \mod.cpu.immdec.imm19_12_20[0] ;
 wire \mod.cpu.immdec.imm19_12_20[1] ;
 wire \mod.cpu.immdec.imm19_12_20[2] ;
 wire \mod.cpu.immdec.imm19_12_20[3] ;
 wire \mod.cpu.immdec.imm19_12_20[5] ;
 wire \mod.cpu.immdec.imm19_12_20[6] ;
 wire \mod.cpu.immdec.imm19_12_20[7] ;
 wire \mod.cpu.immdec.imm19_12_20[8] ;
 wire \mod.cpu.immdec.imm24_20[0] ;
 wire \mod.cpu.immdec.imm24_20[1] ;
 wire \mod.cpu.immdec.imm24_20[2] ;
 wire \mod.cpu.immdec.imm24_20[3] ;
 wire \mod.cpu.immdec.imm24_20[4] ;
 wire \mod.cpu.immdec.imm30_25[0] ;
 wire \mod.cpu.immdec.imm30_25[1] ;
 wire \mod.cpu.immdec.imm30_25[2] ;
 wire \mod.cpu.immdec.imm30_25[3] ;
 wire \mod.cpu.immdec.imm30_25[4] ;
 wire \mod.cpu.immdec.imm30_25[5] ;
 wire \mod.cpu.immdec.imm31 ;
 wire \mod.cpu.immdec.imm7 ;
 wire \mod.cpu.mem_bytecnt[0] ;
 wire \mod.cpu.mem_bytecnt[1] ;
 wire \mod.cpu.mem_if.signbit ;
 wire \mod.cpu.state.ibus_cyc ;
 wire \mod.cpu.state.init_done ;
 wire \mod.cpu.state.o_cnt[2] ;
 wire \mod.cpu.state.o_cnt_r[0] ;
 wire \mod.cpu.state.o_cnt_r[1] ;
 wire \mod.cpu.state.o_cnt_r[2] ;
 wire \mod.cpu.state.o_cnt_r[3] ;
 wire \mod.cpu.state.stage_two_req ;
 wire \mod.u_arbiter.i_wb_cpu_ack ;
 wire \mod.u_scanchain_local.module_data_in[37] ;
 wire \mod.u_scanchain_local.module_data_in[38] ;
 wire \mod.u_scanchain_local.module_data_in[39] ;
 wire \mod.u_scanchain_local.module_data_in[40] ;
 wire \mod.u_scanchain_local.module_data_in[41] ;
 wire \mod.u_scanchain_local.module_data_in[42] ;
 wire \mod.u_scanchain_local.module_data_in[43] ;
 wire \mod.u_scanchain_local.module_data_in[44] ;
 wire \mod.u_scanchain_local.module_data_in[45] ;
 wire \mod.u_scanchain_local.module_data_in[46] ;
 wire \mod.u_scanchain_local.module_data_in[47] ;
 wire \mod.u_scanchain_local.module_data_in[48] ;
 wire \mod.u_scanchain_local.module_data_in[49] ;
 wire \mod.u_scanchain_local.module_data_in[50] ;
 wire \mod.u_scanchain_local.module_data_in[51] ;
 wire \mod.u_scanchain_local.module_data_in[52] ;
 wire \mod.u_scanchain_local.module_data_in[53] ;
 wire \mod.u_scanchain_local.module_data_in[54] ;
 wire \mod.u_scanchain_local.module_data_in[55] ;
 wire \mod.u_scanchain_local.module_data_in[56] ;
 wire \mod.u_scanchain_local.module_data_in[57] ;
 wire \mod.u_scanchain_local.module_data_in[58] ;
 wire \mod.u_scanchain_local.module_data_in[59] ;
 wire \mod.u_scanchain_local.module_data_in[60] ;
 wire \mod.u_scanchain_local.module_data_in[61] ;
 wire \mod.u_scanchain_local.module_data_in[62] ;
 wire \mod.u_scanchain_local.module_data_in[63] ;
 wire \mod.u_scanchain_local.module_data_in[64] ;
 wire \mod.u_scanchain_local.module_data_in[65] ;
 wire \mod.u_scanchain_local.module_data_in[66] ;
 wire \mod.u_scanchain_local.module_data_in[67] ;
 wire \mod.u_scanchain_local.module_data_in[68] ;
 wire \mod.u_scanchain_local.module_data_in[69] ;
 wire \mod.u_scanchain_local.module_data_in[70] ;
 wire \mod.u_scanchain_local.module_data_in[71] ;
 wire \mod.u_scanchain_local.module_data_in[72] ;
 wire \mod.u_scanchain_local.module_data_in[73] ;
 wire \mod.u_scanchain_local.module_data_in[74] ;
 wire \mod.u_scanchain_local.module_data_in[75] ;
 wire \mod.u_scanchain_local.module_data_in[76] ;
 wire \mod.u_scanchain_local.module_data_in[77] ;
 wire \mod.u_scanchain_local.module_data_in[78] ;
 wire \mod.u_scanchain_local.module_data_in[79] ;
 wire \mod.u_scanchain_local.module_data_in[80] ;
 wire \mod.u_scanchain_local.module_data_in[81] ;
 wire \mod.u_scanchain_local.module_data_in[82] ;
 wire \mod.u_scanchain_local.module_data_in[83] ;
 wire \mod.u_scanchain_local.module_data_in[84] ;
 wire \mod.u_scanchain_local.module_data_in[85] ;
 wire \mod.u_scanchain_local.module_data_in[86] ;
 wire \mod.u_scanchain_local.module_data_in[87] ;
 wire \mod.u_scanchain_local.module_data_in[88] ;
 wire \mod.u_scanchain_local.module_data_in[89] ;
 wire \mod.u_scanchain_local.module_data_in[90] ;
 wire \mod.u_scanchain_local.module_data_in[91] ;
 wire \mod.u_scanchain_local.module_data_in[92] ;
 wire \mod.u_scanchain_local.module_data_in[93] ;
 wire \mod.u_scanchain_local.module_data_in[94] ;
 wire \mod.u_scanchain_local.module_data_in[95] ;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net151;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net152;
 wire net180;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;

 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1006_ (.A1(\mod.cpu.state.o_cnt_r[0] ),
    .A2(\mod.cpu.state.o_cnt_r[1] ),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1007_ (.A1(\mod.cpu.state.o_cnt_r[3] ),
    .A2(\mod.cpu.state.o_cnt_r[2] ),
    .A3(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1008_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1009_ (.I(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1010_ (.I(\mod.cpu.decode.co_mem_word ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1011_ (.I(\mod.cpu.bne_or_bge ),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1012_ (.A1(_0606_),
    .A2(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1013_ (.A1(\mod.cpu.bufreg2.i_op_b_sel ),
    .A2(\mod.cpu.bufreg.i_sh_signed ),
    .B(_0608_),
    .C(\mod.cpu.branch_op ),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1014_ (.A1(\mod.cpu.alu.i_rs1 ),
    .A2(\mod.cpu.alu.add_cy_r ),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1015_ (.I(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1016_ (.I(\mod.cpu.bufreg2.i_cnt_done ),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1017_ (.I(\mod.cpu.bufreg2.i_op_b_sel ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1018_ (.A1(\mod.cpu.decode.opcode[0] ),
    .A2(\mod.cpu.decode.opcode[1] ),
    .A3(\mod.cpu.decode.opcode[2] ),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1019_ (.A1(_0613_),
    .A2(\mod.cpu.immdec.imm11_7[0] ),
    .A3(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1020_ (.I(\mod.cpu.decode.opcode[1] ),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1021_ (.A1(\mod.cpu.decode.opcode[0] ),
    .A2(_0616_),
    .A3(\mod.cpu.decode.opcode[2] ),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1022_ (.A1(\mod.cpu.bufreg2.i_op_b_sel ),
    .A2(_0617_),
    .B(\mod.cpu.immdec.imm24_20[0] ),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1023_ (.I(\mod.cpu.decode.opcode[2] ),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1024_ (.A1(_0619_),
    .A2(\mod.cpu.branch_op ),
    .A3(\mod.cpu.csr_d_sel ),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1025_ (.A1(\mod.cpu.bufreg2.i_cnt_done ),
    .A2(\mod.cpu.immdec.imm31 ),
    .A3(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1026_ (.A1(_0612_),
    .A2(_0615_),
    .A3(_0618_),
    .B(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1027_ (.I0(\mod.cpu.bufreg2.i_rs2 ),
    .I1(_0622_),
    .S(_0613_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1028_ (.A1(_0609_),
    .A2(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1029_ (.I(\mod.cpu.alu.i_rs1 ),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1030_ (.A1(_0625_),
    .A2(\mod.cpu.alu.add_cy_r ),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1031_ (.A1(_0611_),
    .A2(_0624_),
    .B(_0626_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1032_ (.A1(_0605_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1033_ (.A1(_0605_),
    .A2(_0609_),
    .B(_0628_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1034_ (.I(net2),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1035_ (.I(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1036_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1037_ (.I0(net1),
    .I1(\mod.cpu.immdec.imm24_20[0] ),
    .S(_0631_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1038_ (.I(_0632_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1039_ (.I0(\mod.cpu.bufreg2.i_rs2 ),
    .I1(\mod.cpu.immdec.imm24_20[1] ),
    .S(_0631_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1040_ (.I(_0633_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1041_ (.I(_0625_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1042_ (.I0(_0634_),
    .I1(\mod.cpu.immdec.imm24_20[2] ),
    .S(_0631_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1043_ (.I(_0635_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1044_ (.I0(\mod.cpu.i_rf_ready ),
    .I1(\mod.cpu.immdec.imm24_20[3] ),
    .S(_0631_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1045_ (.I(_0636_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1046_ (.I(_0630_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1047_ (.I0(\mod.cpu.i_timer_irq ),
    .I1(\mod.cpu.immdec.imm24_20[4] ),
    .S(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1048_ (.I(_0638_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1049_ (.I(\mod.u_arbiter.i_wb_cpu_ack ),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1050_ (.I0(_0639_),
    .I1(\mod.cpu.csr_imm ),
    .S(_0637_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1051_ (.I(_0640_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1052_ (.I0(\mod.cpu.bufreg2.i_dat[0] ),
    .I1(\mod.cpu.immdec.imm19_12_20[5] ),
    .S(_0637_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1053_ (.I(_0641_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1054_ (.I0(\mod.cpu.bufreg2.i_dat[1] ),
    .I1(\mod.cpu.immdec.imm19_12_20[6] ),
    .S(_0637_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1055_ (.I(_0642_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1056_ (.I(_0630_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1057_ (.I0(\mod.cpu.bufreg2.i_dat[2] ),
    .I1(\mod.cpu.immdec.imm19_12_20[7] ),
    .S(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1058_ (.I(_0644_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1059_ (.I(\mod.cpu.immdec.imm19_12_20[8] ),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1060_ (.I(net2),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1061_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1062_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1063_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1064_ (.I(_0646_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1065_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1066_ (.I(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1067_ (.A1(\mod.cpu.bufreg2.i_dat[3] ),
    .A2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1068_ (.A1(_0645_),
    .A2(_0649_),
    .B(_0653_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1069_ (.I(\mod.cpu.bufreg2.i_dat[5] ),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1070_ (.I(_0619_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1071_ (.I(\mod.cpu.csr_d_sel ),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1072_ (.I(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1073_ (.I(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1074_ (.A1(_0610_),
    .A2(_0624_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1075_ (.A1(_0658_),
    .A2(_0608_),
    .A3(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1076_ (.I(_0606_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1077_ (.A1(\mod.cpu.mem_bytecnt[0] ),
    .A2(\mod.cpu.state.o_cnt[2] ),
    .A3(\mod.cpu.mem_bytecnt[1] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1078_ (.A1(\mod.cpu.state.o_cnt_r[0] ),
    .A2(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1079_ (.A1(_0657_),
    .A2(_0661_),
    .A3(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1080_ (.I(_0623_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1081_ (.A1(_0661_),
    .A2(_0634_),
    .A3(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1082_ (.I(\mod.cpu.bne_or_bge ),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1083_ (.A1(_0625_),
    .A2(_0665_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1084_ (.A1(_0667_),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1085_ (.A1(_0625_),
    .A2(_0665_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1086_ (.A1(_0657_),
    .A2(_0666_),
    .A3(_0669_),
    .A4(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1087_ (.A1(_0656_),
    .A2(\mod.cpu.bufreg2.dat[5] ),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1088_ (.I(\mod.cpu.state.init_done ),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1089_ (.I(_0619_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1090_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1091_ (.I(\mod.cpu.decode.co_mem_word ),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1092_ (.A1(_0675_),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1093_ (.A1(_0673_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1094_ (.I(\mod.cpu.state.o_cnt_r[3] ),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1095_ (.I(\mod.cpu.state.o_cnt_r[2] ),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1096_ (.A1(_0679_),
    .A2(_0680_),
    .A3(_0602_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1097_ (.I(_0674_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1098_ (.I(\mod.cpu.branch_op ),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1099_ (.I(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1100_ (.A1(\mod.cpu.decode.co_mem_word ),
    .A2(\mod.cpu.bne_or_bge ),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1101_ (.I(\mod.cpu.decode.opcode[0] ),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1102_ (.A1(_0686_),
    .A2(\mod.cpu.branch_op ),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1103_ (.A1(\mod.cpu.csr_d_sel ),
    .A2(\mod.cpu.decode.co_mem_word ),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1104_ (.A1(_0685_),
    .A2(_0687_),
    .A3(_0688_),
    .B(_0619_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1105_ (.I(\mod.cpu.state.init_done ),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1106_ (.A1(_0682_),
    .A2(_0684_),
    .B1(_0689_),
    .B2(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1107_ (.A1(\mod.cpu.state.stage_two_req ),
    .A2(_0672_),
    .A3(_0678_),
    .B1(_0681_),
    .B2(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1108_ (.A1(\mod.cpu.bufreg.lsb[0] ),
    .A2(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1109_ (.A1(\mod.cpu.alu.cmp_r ),
    .A2(_0664_),
    .B(_0671_),
    .C(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1110_ (.A1(_0660_),
    .A2(_0694_),
    .B(_0687_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1111_ (.A1(_0655_),
    .A2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1112_ (.I(\mod.cpu.decode.opcode[0] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1113_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1114_ (.I(_0675_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1115_ (.A1(_0698_),
    .A2(_0699_),
    .A3(_0684_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1116_ (.I(_0683_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1117_ (.A1(_0675_),
    .A2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1118_ (.I(\mod.cpu.bufreg2.i_op_b_sel ),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1119_ (.A1(_0683_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1120_ (.A1(_0686_),
    .A2(_0616_),
    .B1(\mod.cpu.decode.co_ebreak ),
    .B2(_0702_),
    .C(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1121_ (.A1(_0614_),
    .A2(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1122_ (.A1(\mod.cpu.ctrl.o_ibus_adr[0] ),
    .A2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1123_ (.A1(\mod.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_0707_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1124_ (.I(\mod.cpu.mem_bytecnt[1] ),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1125_ (.A1(\mod.cpu.mem_bytecnt[0] ),
    .A2(\mod.cpu.state.o_cnt[2] ),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1126_ (.A1(_0709_),
    .A2(_0710_),
    .B(_0622_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1127_ (.A1(_0700_),
    .A2(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1128_ (.A1(_0693_),
    .A2(_0700_),
    .B(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1129_ (.A1(_0708_),
    .A2(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1130_ (.A1(_0708_),
    .A2(_0713_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1131_ (.A1(_0663_),
    .A2(_0714_),
    .A3(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1132_ (.I(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1133_ (.I(_0676_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1134_ (.I(\mod.cpu.mem_if.signbit ),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1135_ (.I(\mod.cpu.mem_bytecnt[0] ),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1136_ (.A1(_0607_),
    .A2(_0720_),
    .B(_0709_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1137_ (.I(\mod.cpu.bufreg.lsb[1] ),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1138_ (.I0(\mod.cpu.bufreg2.dat[0] ),
    .I1(\mod.cpu.bufreg2.dat[8] ),
    .I2(\mod.cpu.bufreg2.dat[16] ),
    .I3(\mod.cpu.bufreg2.dat[24] ),
    .S0(\mod.cpu.bufreg.lsb[0] ),
    .S1(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1139_ (.A1(_0718_),
    .A2(_0721_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1140_ (.A1(_0718_),
    .A2(_0719_),
    .A3(_0721_),
    .B(_0724_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1141_ (.I(_0686_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1142_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1143_ (.A1(_0658_),
    .A2(_0724_),
    .B(_0726_),
    .C(_0655_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1144_ (.I(_0629_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1145_ (.I(_0683_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1146_ (.I(_0662_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1147_ (.A1(_0680_),
    .A2(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1148_ (.A1(\mod.cpu.ctrl.pc_plus_4_cy_r ),
    .A2(\mod.cpu.ctrl.o_ibus_adr[0] ),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1149_ (.A1(_0731_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1150_ (.A1(_0726_),
    .A2(_0729_),
    .A3(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1151_ (.A1(_0728_),
    .A2(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1152_ (.A1(_0700_),
    .A2(_0717_),
    .B1(_0101_),
    .B2(_0727_),
    .C(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1153_ (.A1(_0654_),
    .A2(_0649_),
    .B1(_0696_),
    .B2(_0736_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1154_ (.I(\mod.cpu.bufreg2.i_dat[7] ),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1155_ (.I(_0728_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1156_ (.A1(_0690_),
    .A2(_0689_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1157_ (.A1(_0603_),
    .A2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1158_ (.A1(\mod.cpu.immdec.imm11_7[1] ),
    .A2(\mod.cpu.immdec.imm11_7[2] ),
    .A3(\mod.cpu.immdec.imm11_7[3] ),
    .A4(\mod.cpu.immdec.imm11_7[0] ),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1159_ (.A1(_0686_),
    .A2(_0684_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1160_ (.A1(_0725_),
    .A2(_0703_),
    .B(_0742_),
    .C(_0682_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1161_ (.A1(\mod.cpu.immdec.imm11_7[4] ),
    .A2(_0741_),
    .B(_0743_),
    .C(_0728_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1162_ (.A1(_0737_),
    .A2(_0738_),
    .B1(_0740_),
    .B2(_0744_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1163_ (.I0(\mod.cpu.bufreg2.i_dat[13] ),
    .I1(\mod.cpu.immdec.imm11_7[0] ),
    .S(_0643_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1164_ (.I(_0745_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1165_ (.I0(\mod.cpu.bufreg2.i_dat[14] ),
    .I1(\mod.cpu.immdec.imm11_7[1] ),
    .S(_0643_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1166_ (.I(_0746_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1167_ (.I(\mod.cpu.immdec.imm11_7[2] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1168_ (.I(_0648_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1169_ (.I(_0651_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1170_ (.A1(\mod.cpu.bufreg2.i_dat[15] ),
    .A2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1171_ (.A1(_0747_),
    .A2(_0748_),
    .B(_0750_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1172_ (.I(\mod.cpu.immdec.imm11_7[3] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1173_ (.A1(\mod.cpu.bufreg2.i_dat[16] ),
    .A2(_0749_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1174_ (.A1(_0751_),
    .A2(_0748_),
    .B(_0752_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1175_ (.I0(\mod.cpu.bufreg2.i_dat[17] ),
    .I1(\mod.cpu.immdec.imm11_7[4] ),
    .S(_0643_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1176_ (.I(_0753_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1177_ (.I(_0650_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1178_ (.I(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1179_ (.I(net3),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1180_ (.A1(_0756_),
    .A2(\mod.cpu.state.ibus_cyc ),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1181_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1182_ (.I(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1183_ (.I(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1184_ (.I(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1185_ (.I(_0761_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1186_ (.A1(\mod.cpu.bufreg2.i_dat[18] ),
    .A2(_0749_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1187_ (.A1(_0755_),
    .A2(_0762_),
    .B(_0763_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1188_ (.I(_0739_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1189_ (.A1(_0612_),
    .A2(_0764_),
    .B(_0677_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1190_ (.I(\mod.cpu.bufreg2.dat[5] ),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1191_ (.A1(\mod.cpu.bufreg2.dat[0] ),
    .A2(\mod.cpu.bufreg2.dat[1] ),
    .A3(\mod.cpu.bufreg2.dat[2] ),
    .A4(\mod.cpu.bufreg2.dat[3] ),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1192_ (.A1(\mod.cpu.bufreg2.dat[4] ),
    .A2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1193_ (.A1(_0766_),
    .A2(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1194_ (.A1(_0739_),
    .A2(_0677_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1195_ (.I(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1196_ (.A1(\mod.cpu.bufreg2.dat[6] ),
    .A2(_0765_),
    .B1(_0769_),
    .B2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1197_ (.A1(_0658_),
    .A2(_0661_),
    .A3(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1198_ (.A1(_0756_),
    .A2(\mod.cpu.state.ibus_cyc ),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1199_ (.A1(_0639_),
    .A2(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1200_ (.I(_0775_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1201_ (.I(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1202_ (.I(_0729_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1203_ (.A1(_0655_),
    .A2(_0773_),
    .B(_0777_),
    .C(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1204_ (.I(_0629_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1205_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1206_ (.I(_0681_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1207_ (.I(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1208_ (.A1(_0673_),
    .A2(_0781_),
    .A3(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1209_ (.A1(\mod.cpu.bufreg2.i_dat[19] ),
    .A2(_0749_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1210_ (.A1(_0779_),
    .A2(_0784_),
    .B(_0785_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1211_ (.A1(_0673_),
    .A2(_0701_),
    .A3(_0783_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1212_ (.I(_0774_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1213_ (.I(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1214_ (.A1(_0655_),
    .A2(_0786_),
    .B(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1215_ (.I(_0630_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1216_ (.I0(\mod.cpu.bufreg2.i_dat[20] ),
    .I1(_0789_),
    .S(_0790_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1217_ (.I(_0791_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1218_ (.I(\mod.cpu.bufreg2.i_dat[21] ),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1219_ (.I(_0780_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1220_ (.I(_0774_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1221_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1222_ (.A1(_0703_),
    .A2(_0793_),
    .A3(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1223_ (.A1(_0792_),
    .A2(_0738_),
    .B(_0796_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1224_ (.I(\mod.cpu.bufreg.lsb[0] ),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1225_ (.A1(_0797_),
    .A2(_0722_),
    .B(_0728_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1226_ (.A1(\mod.cpu.bufreg2.i_dat[22] ),
    .A2(_0738_),
    .B(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1227_ (.I(_0799_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1228_ (.A1(_0667_),
    .A2(_0797_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1229_ (.A1(_0718_),
    .A2(_0651_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1230_ (.A1(_0722_),
    .A2(_0800_),
    .B(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1231_ (.A1(\mod.cpu.bufreg2.i_dat[23] ),
    .A2(_0793_),
    .B(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1232_ (.I(_0803_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1233_ (.I(\mod.cpu.bufreg2.i_dat[24] ),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1234_ (.I(_0797_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1235_ (.I(_0722_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1236_ (.A1(_0805_),
    .A2(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1237_ (.A1(_0804_),
    .A2(_0649_),
    .B1(_0807_),
    .B2(_0801_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1238_ (.I(\mod.cpu.bufreg2.i_dat[25] ),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1239_ (.A1(_0667_),
    .A2(_0797_),
    .B(_0806_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1240_ (.A1(_0808_),
    .A2(_0649_),
    .B1(_0801_),
    .B2(_0809_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1241_ (.I(\mod.cpu.bufreg2.dat[0] ),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1242_ (.I0(\mod.cpu.bufreg2.i_dat[26] ),
    .I1(_0810_),
    .S(_0790_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1243_ (.I(_0811_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1244_ (.I(\mod.cpu.bufreg2.dat[1] ),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1245_ (.I0(\mod.cpu.bufreg2.i_dat[27] ),
    .I1(_0812_),
    .S(_0790_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1246_ (.I(_0813_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1247_ (.I(\mod.cpu.bufreg2.dat[2] ),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1248_ (.I0(\mod.cpu.bufreg2.i_dat[28] ),
    .I1(_0814_),
    .S(_0790_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1249_ (.I(_0815_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1250_ (.I(_0629_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1251_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1252_ (.I0(\mod.cpu.bufreg2.i_dat[29] ),
    .I1(\mod.cpu.bufreg2.dat[3] ),
    .S(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1253_ (.I(_0818_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1254_ (.I(\mod.cpu.bufreg2.dat[4] ),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1255_ (.I0(\mod.cpu.bufreg2.i_dat[30] ),
    .I1(_0819_),
    .S(_0817_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1256_ (.I(_0820_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1257_ (.I0(\mod.cpu.bufreg2.i_dat[31] ),
    .I1(_0766_),
    .S(_0817_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1258_ (.I(_0821_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1259_ (.I0(\mod.u_scanchain_local.module_data_in[37] ),
    .I1(\mod.cpu.bufreg2.dat[6] ),
    .S(_0817_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1260_ (.I(_0822_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1261_ (.I(_0816_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1262_ (.I0(\mod.u_scanchain_local.module_data_in[38] ),
    .I1(\mod.cpu.bufreg2.dat[7] ),
    .S(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1263_ (.I(_0824_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1264_ (.I0(\mod.u_scanchain_local.module_data_in[39] ),
    .I1(\mod.cpu.bufreg2.dat[8] ),
    .S(_0823_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1265_ (.I(_0825_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1266_ (.I0(\mod.u_scanchain_local.module_data_in[40] ),
    .I1(\mod.cpu.bufreg2.dat[9] ),
    .S(_0823_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1267_ (.I(_0826_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1268_ (.I0(\mod.u_scanchain_local.module_data_in[41] ),
    .I1(\mod.cpu.bufreg2.dat[10] ),
    .S(_0823_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1269_ (.I(_0827_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1270_ (.I(_0816_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1271_ (.I0(\mod.u_scanchain_local.module_data_in[42] ),
    .I1(\mod.cpu.bufreg2.dat[11] ),
    .S(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1272_ (.I(_0829_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1273_ (.I0(\mod.u_scanchain_local.module_data_in[43] ),
    .I1(\mod.cpu.bufreg2.dat[12] ),
    .S(_0828_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1274_ (.I(_0830_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1275_ (.I0(\mod.u_scanchain_local.module_data_in[44] ),
    .I1(\mod.cpu.bufreg2.dat[13] ),
    .S(_0828_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1276_ (.I(_0831_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1277_ (.I0(\mod.u_scanchain_local.module_data_in[45] ),
    .I1(\mod.cpu.bufreg2.dat[14] ),
    .S(_0828_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1278_ (.I(_0832_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1279_ (.I(_0816_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1280_ (.I0(\mod.u_scanchain_local.module_data_in[46] ),
    .I1(\mod.cpu.bufreg2.dat[15] ),
    .S(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1281_ (.I(_0834_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1282_ (.I0(\mod.u_scanchain_local.module_data_in[47] ),
    .I1(\mod.cpu.bufreg2.dat[16] ),
    .S(_0833_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1283_ (.I(_0835_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1284_ (.I0(\mod.u_scanchain_local.module_data_in[48] ),
    .I1(\mod.cpu.bufreg2.dat[17] ),
    .S(_0833_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1285_ (.I(_0836_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1286_ (.I0(\mod.u_scanchain_local.module_data_in[49] ),
    .I1(\mod.cpu.bufreg2.dat[18] ),
    .S(_0833_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1287_ (.I(_0837_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1288_ (.I(_0780_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1289_ (.I0(\mod.u_scanchain_local.module_data_in[50] ),
    .I1(\mod.cpu.bufreg2.dat[19] ),
    .S(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1290_ (.I(_0839_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1291_ (.I0(\mod.u_scanchain_local.module_data_in[51] ),
    .I1(\mod.cpu.bufreg2.dat[20] ),
    .S(_0838_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1292_ (.I(_0840_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1293_ (.I0(\mod.u_scanchain_local.module_data_in[52] ),
    .I1(\mod.cpu.bufreg2.dat[21] ),
    .S(_0838_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1294_ (.I(_0841_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1295_ (.I0(\mod.u_scanchain_local.module_data_in[53] ),
    .I1(\mod.cpu.bufreg2.dat[22] ),
    .S(_0838_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1296_ (.I(_0842_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1297_ (.I(_0780_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1298_ (.I0(\mod.u_scanchain_local.module_data_in[54] ),
    .I1(\mod.cpu.bufreg2.dat[23] ),
    .S(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1299_ (.I(_0844_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1300_ (.I0(\mod.u_scanchain_local.module_data_in[55] ),
    .I1(\mod.cpu.bufreg2.dat[24] ),
    .S(_0843_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1301_ (.I(_0845_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1302_ (.I0(\mod.u_scanchain_local.module_data_in[56] ),
    .I1(\mod.cpu.bufreg2.dat[25] ),
    .S(_0843_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1303_ (.I(_0846_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1304_ (.I(\mod.cpu.bufreg2.dat[26] ),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1305_ (.A1(_0652_),
    .A2(\mod.u_scanchain_local.module_data_in[57] ),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1306_ (.A1(_0847_),
    .A2(_0748_),
    .B(_0848_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1307_ (.I0(\mod.u_scanchain_local.module_data_in[58] ),
    .I1(\mod.cpu.bufreg2.dat[27] ),
    .S(_0843_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1308_ (.I(_0849_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1309_ (.I0(\mod.u_scanchain_local.module_data_in[59] ),
    .I1(\mod.cpu.bufreg2.dat[28] ),
    .S(_0781_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1310_ (.I(_0850_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1311_ (.I0(\mod.u_scanchain_local.module_data_in[60] ),
    .I1(\mod.cpu.bufreg2.dat[29] ),
    .S(_0781_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1312_ (.I(_0851_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1313_ (.I(\mod.cpu.bufreg2.dat[30] ),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1314_ (.A1(_0652_),
    .A2(\mod.u_scanchain_local.module_data_in[61] ),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1315_ (.A1(_0852_),
    .A2(_0748_),
    .B(_0853_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1316_ (.I(\mod.cpu.bufreg2.dat[31] ),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1317_ (.I(_0754_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1318_ (.A1(_0652_),
    .A2(\mod.u_scanchain_local.module_data_in[62] ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1319_ (.A1(_0854_),
    .A2(_0855_),
    .B(_0856_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1320_ (.I(_0651_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1321_ (.A1(_0857_),
    .A2(\mod.u_scanchain_local.module_data_in[63] ),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1322_ (.I(\mod.cpu.ctrl.o_ibus_adr[0] ),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1323_ (.I(_0757_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1324_ (.I(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1325_ (.A1(_0859_),
    .A2(_0793_),
    .A3(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1326_ (.A1(_0858_),
    .A2(_0862_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1327_ (.A1(_0857_),
    .A2(\mod.u_scanchain_local.module_data_in[64] ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1328_ (.A1(\mod.cpu.ctrl.o_ibus_adr[1] ),
    .A2(_0793_),
    .A3(_0861_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1329_ (.A1(_0863_),
    .A2(_0864_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1330_ (.I(\mod.u_scanchain_local.module_data_in[65] ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1331_ (.A1(\mod.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_0861_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1332_ (.I(_0650_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1333_ (.I(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1334_ (.A1(\mod.cpu.bufreg.data[2] ),
    .A2(_0795_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1335_ (.A1(_0855_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0869_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1336_ (.I(\mod.u_scanchain_local.module_data_in[66] ),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1337_ (.A1(\mod.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0861_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1338_ (.A1(\mod.cpu.bufreg.data[3] ),
    .A2(_0795_),
    .B(_0868_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1339_ (.A1(_0855_),
    .A2(_0870_),
    .B1(_0871_),
    .B2(_0872_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1340_ (.I(\mod.u_scanchain_local.module_data_in[67] ),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1341_ (.I(_0860_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1342_ (.A1(\mod.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1343_ (.A1(\mod.cpu.bufreg.data[4] ),
    .A2(_0795_),
    .B(_0868_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1344_ (.A1(_0855_),
    .A2(_0873_),
    .B1(_0875_),
    .B2(_0876_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1345_ (.I(_0650_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1346_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1347_ (.I(\mod.u_scanchain_local.module_data_in[68] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1348_ (.A1(\mod.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_0874_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1349_ (.I(_0794_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1350_ (.A1(\mod.cpu.bufreg.data[5] ),
    .A2(_0881_),
    .B(_0868_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1351_ (.A1(_0878_),
    .A2(_0879_),
    .B1(_0880_),
    .B2(_0882_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1352_ (.I(\mod.u_scanchain_local.module_data_in[69] ),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1353_ (.A1(\mod.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_0874_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1354_ (.I(_0867_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1355_ (.A1(\mod.cpu.bufreg.data[6] ),
    .A2(_0881_),
    .B(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1356_ (.A1(_0878_),
    .A2(_0883_),
    .B1(_0884_),
    .B2(_0886_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1357_ (.I(\mod.u_scanchain_local.module_data_in[70] ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1358_ (.A1(\mod.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0874_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1359_ (.A1(\mod.cpu.bufreg.data[7] ),
    .A2(_0881_),
    .B(_0885_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1360_ (.A1(_0878_),
    .A2(_0887_),
    .B1(_0888_),
    .B2(_0889_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1361_ (.I(\mod.u_scanchain_local.module_data_in[71] ),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1362_ (.I(_0860_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1363_ (.A1(\mod.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1364_ (.A1(\mod.cpu.bufreg.data[8] ),
    .A2(_0881_),
    .B(_0885_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1365_ (.A1(_0878_),
    .A2(_0890_),
    .B1(_0892_),
    .B2(_0893_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1366_ (.I(_0877_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1367_ (.I(\mod.u_scanchain_local.module_data_in[72] ),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1368_ (.A1(\mod.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0891_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1369_ (.I(_0794_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1370_ (.A1(\mod.cpu.bufreg.data[9] ),
    .A2(_0897_),
    .B(_0885_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1371_ (.A1(_0894_),
    .A2(_0895_),
    .B1(_0896_),
    .B2(_0898_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1372_ (.I(\mod.u_scanchain_local.module_data_in[73] ),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1373_ (.A1(\mod.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0891_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1374_ (.I(_0867_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1375_ (.A1(\mod.cpu.bufreg.data[10] ),
    .A2(_0897_),
    .B(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1376_ (.A1(_0894_),
    .A2(_0899_),
    .B1(_0900_),
    .B2(_0902_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1377_ (.I(\mod.u_scanchain_local.module_data_in[74] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1378_ (.A1(\mod.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_0891_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1379_ (.A1(\mod.cpu.bufreg.data[11] ),
    .A2(_0897_),
    .B(_0901_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1380_ (.A1(_0894_),
    .A2(_0903_),
    .B1(_0904_),
    .B2(_0905_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1381_ (.I(\mod.u_scanchain_local.module_data_in[75] ),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1382_ (.I(_0860_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1383_ (.A1(\mod.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1384_ (.A1(\mod.cpu.bufreg.data[12] ),
    .A2(_0897_),
    .B(_0901_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1385_ (.A1(_0894_),
    .A2(_0906_),
    .B1(_0908_),
    .B2(_0909_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1386_ (.I(_0877_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1387_ (.I(\mod.u_scanchain_local.module_data_in[76] ),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1388_ (.A1(\mod.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_0907_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1389_ (.I(_0794_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1390_ (.A1(\mod.cpu.bufreg.data[13] ),
    .A2(_0913_),
    .B(_0901_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1391_ (.A1(_0910_),
    .A2(_0911_),
    .B1(_0912_),
    .B2(_0914_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1392_ (.I(\mod.u_scanchain_local.module_data_in[77] ),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1393_ (.A1(\mod.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0907_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1394_ (.I(_0867_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1395_ (.A1(\mod.cpu.bufreg.data[14] ),
    .A2(_0913_),
    .B(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1396_ (.A1(_0910_),
    .A2(_0915_),
    .B1(_0916_),
    .B2(_0918_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1397_ (.I(\mod.u_scanchain_local.module_data_in[78] ),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1398_ (.A1(\mod.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_0907_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1399_ (.A1(\mod.cpu.bufreg.data[15] ),
    .A2(_0913_),
    .B(_0917_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1400_ (.A1(_0910_),
    .A2(_0919_),
    .B1(_0920_),
    .B2(_0921_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1401_ (.I(\mod.u_scanchain_local.module_data_in[79] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1402_ (.I(_0757_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1403_ (.I(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1404_ (.A1(\mod.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1405_ (.A1(\mod.cpu.bufreg.data[16] ),
    .A2(_0913_),
    .B(_0917_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1406_ (.A1(_0910_),
    .A2(_0922_),
    .B1(_0925_),
    .B2(_0926_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1407_ (.I(_0877_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1408_ (.I(\mod.u_scanchain_local.module_data_in[80] ),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1409_ (.A1(\mod.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_0924_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1410_ (.I(_0787_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1411_ (.A1(\mod.cpu.bufreg.data[17] ),
    .A2(_0930_),
    .B(_0917_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1412_ (.A1(_0927_),
    .A2(_0928_),
    .B1(_0929_),
    .B2(_0931_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1413_ (.I(\mod.u_scanchain_local.module_data_in[81] ),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1414_ (.A1(\mod.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0924_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1415_ (.I(_0647_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1416_ (.A1(\mod.cpu.bufreg.data[18] ),
    .A2(_0930_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1417_ (.A1(_0927_),
    .A2(_0932_),
    .B1(_0933_),
    .B2(_0935_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1418_ (.I(\mod.u_scanchain_local.module_data_in[82] ),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1419_ (.A1(\mod.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_0924_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1420_ (.A1(\mod.cpu.bufreg.data[19] ),
    .A2(_0930_),
    .B(_0934_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1421_ (.A1(_0927_),
    .A2(_0936_),
    .B1(_0937_),
    .B2(_0938_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1422_ (.I(\mod.u_scanchain_local.module_data_in[83] ),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1423_ (.I(_0923_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1424_ (.A1(\mod.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1425_ (.A1(\mod.cpu.bufreg.data[20] ),
    .A2(_0930_),
    .B(_0934_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1426_ (.A1(_0927_),
    .A2(_0939_),
    .B1(_0941_),
    .B2(_0942_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1427_ (.I(_0754_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1428_ (.I(\mod.u_scanchain_local.module_data_in[84] ),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1429_ (.A1(\mod.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0940_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1430_ (.I(_0787_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1431_ (.A1(\mod.cpu.bufreg.data[21] ),
    .A2(_0946_),
    .B(_0934_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1432_ (.A1(_0943_),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0947_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1433_ (.I(\mod.u_scanchain_local.module_data_in[85] ),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1434_ (.A1(\mod.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0940_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1435_ (.I(_0647_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1436_ (.A1(\mod.cpu.bufreg.data[22] ),
    .A2(_0946_),
    .B(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1437_ (.A1(_0943_),
    .A2(_0948_),
    .B1(_0949_),
    .B2(_0951_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1438_ (.I(\mod.u_scanchain_local.module_data_in[86] ),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1439_ (.A1(\mod.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0940_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1440_ (.A1(\mod.cpu.bufreg.data[23] ),
    .A2(_0946_),
    .B(_0950_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1441_ (.A1(_0943_),
    .A2(_0952_),
    .B1(_0953_),
    .B2(_0954_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1442_ (.I(\mod.u_scanchain_local.module_data_in[87] ),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1443_ (.I(_0923_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1444_ (.A1(\mod.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1445_ (.A1(\mod.cpu.bufreg.data[24] ),
    .A2(_0946_),
    .B(_0950_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1446_ (.A1(_0943_),
    .A2(_0955_),
    .B1(_0957_),
    .B2(_0958_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1447_ (.I(_0754_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1448_ (.I(\mod.u_scanchain_local.module_data_in[88] ),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1449_ (.A1(\mod.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0956_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1450_ (.I(_0787_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1451_ (.A1(\mod.cpu.bufreg.data[25] ),
    .A2(_0962_),
    .B(_0950_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1452_ (.A1(_0959_),
    .A2(_0960_),
    .B1(_0961_),
    .B2(_0963_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1453_ (.I(\mod.u_scanchain_local.module_data_in[89] ),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1454_ (.A1(\mod.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0956_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1455_ (.I(_0647_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1456_ (.A1(\mod.cpu.bufreg.data[26] ),
    .A2(_0962_),
    .B(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1457_ (.A1(_0959_),
    .A2(_0964_),
    .B1(_0965_),
    .B2(_0967_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1458_ (.I(\mod.u_scanchain_local.module_data_in[90] ),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1459_ (.A1(\mod.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_0956_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1460_ (.A1(\mod.cpu.bufreg.data[27] ),
    .A2(_0962_),
    .B(_0966_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1461_ (.A1(_0959_),
    .A2(_0968_),
    .B1(_0969_),
    .B2(_0970_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1462_ (.I(\mod.u_scanchain_local.module_data_in[91] ),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1463_ (.I(_0923_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1464_ (.A1(\mod.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1465_ (.A1(\mod.cpu.bufreg.data[28] ),
    .A2(_0962_),
    .B(_0966_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1466_ (.A1(_0959_),
    .A2(_0971_),
    .B1(_0973_),
    .B2(_0974_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1467_ (.I(\mod.u_scanchain_local.module_data_in[92] ),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1468_ (.A1(\mod.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0972_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1469_ (.A1(\mod.cpu.bufreg.data[29] ),
    .A2(_0788_),
    .B(_0966_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1470_ (.A1(_0755_),
    .A2(_0975_),
    .B1(_0976_),
    .B2(_0977_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1471_ (.I(\mod.u_scanchain_local.module_data_in[93] ),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1472_ (.A1(\mod.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_0972_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1473_ (.A1(\mod.cpu.bufreg.data[30] ),
    .A2(_0788_),
    .B(_0648_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1474_ (.A1(_0755_),
    .A2(_0978_),
    .B1(_0979_),
    .B2(_0980_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1475_ (.I(\mod.u_scanchain_local.module_data_in[94] ),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1476_ (.A1(\mod.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0972_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1477_ (.A1(\mod.cpu.bufreg.data[31] ),
    .A2(_0788_),
    .B(_0648_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1478_ (.A1(_0755_),
    .A2(_0981_),
    .B1(_0982_),
    .B2(_0983_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1479_ (.I(_0616_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1480_ (.A1(_0984_),
    .A2(_0729_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1481_ (.A1(_0698_),
    .A2(_0684_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1482_ (.A1(_0634_),
    .A2(\mod.cpu.bufreg.c_r ),
    .A3(_0985_),
    .A4(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1483_ (.A1(_0634_),
    .A2(_0985_),
    .A3(_0986_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1484_ (.A1(\mod.cpu.bufreg.c_r ),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1485_ (.A1(_0725_),
    .A2(_0616_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1486_ (.A1(_0701_),
    .A2(_0663_),
    .A3(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1487_ (.A1(_0699_),
    .A2(_0622_),
    .A3(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1488_ (.A1(_0989_),
    .A2(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1489_ (.A1(_0782_),
    .A2(_0691_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1490_ (.A1(\mod.cpu.state.stage_two_req ),
    .A2(_0672_),
    .A3(_0678_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1491_ (.A1(_0994_),
    .A2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1492_ (.A1(_0987_),
    .A2(_0993_),
    .B(_0996_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1493_ (.A1(_0859_),
    .A2(\mod.cpu.ctrl.pc_plus_offset_cy_r ),
    .A3(_0706_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1494_ (.A1(_0997_),
    .A2(_0714_),
    .B(_0740_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1495_ (.A1(\mod.cpu.ctrl.pc_plus_4_cy_r ),
    .A2(_0859_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1496_ (.A1(_0680_),
    .A2(_0730_),
    .A3(_0732_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1497_ (.A1(_0998_),
    .A2(_0999_),
    .B(_0740_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1498_ (.A1(\mod.cpu.bufreg2.i_dat[4] ),
    .A2(_0857_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1499_ (.I(_1000_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1500_ (.I(\mod.cpu.bufreg2.i_dat[6] ),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1501_ (.I(_0781_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1502_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1503_ (.I(\mod.cpu.bufreg2.i_dat[8] ),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1504_ (.A1(_1003_),
    .A2(_1002_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1505_ (.I(\mod.cpu.bufreg2.i_dat[9] ),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1506_ (.A1(_1004_),
    .A2(_1002_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1507_ (.I(\mod.cpu.bufreg2.i_dat[10] ),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1508_ (.A1(_1005_),
    .A2(_1002_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1509_ (.I(\mod.cpu.bufreg2.i_dat[11] ),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1510_ (.A1(_0247_),
    .A2(_0738_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1511_ (.A1(\mod.cpu.bufreg2.i_dat[12] ),
    .A2(_0857_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1512_ (.I(_0248_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1513_ (.I(net3),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1514_ (.A1(_0604_),
    .A2(_0739_),
    .B(_0249_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1515_ (.I(_0250_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1516_ (.I(_0760_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1517_ (.I(_0249_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1518_ (.A1(_0253_),
    .A2(_0612_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1519_ (.A1(_0252_),
    .A2(_0254_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1520_ (.A1(\mod.cpu.state.ibus_cyc ),
    .A2(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1521_ (.A1(_0251_),
    .A2(_0255_),
    .B(_0256_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1522_ (.A1(\mod.cpu.ctrl.i_jump ),
    .A2(_0254_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1523_ (.A1(\mod.cpu.state.o_cnt_r[0] ),
    .A2(_0730_),
    .B(\mod.cpu.alu.cmp_r ),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1524_ (.A1(_0657_),
    .A2(_0718_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1525_ (.A1(_0659_),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1526_ (.A1(_0656_),
    .A2(\mod.cpu.bne_or_bge ),
    .B(_0676_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1527_ (.A1(_0668_),
    .A2(_0670_),
    .A3(_0261_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1528_ (.A1(_0627_),
    .A2(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1529_ (.A1(_0258_),
    .A2(_0260_),
    .B1(_0263_),
    .B2(_0259_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1530_ (.A1(_0667_),
    .A2(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1531_ (.I(_0612_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1532_ (.A1(_0249_),
    .A2(_0266_),
    .A3(_0764_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1533_ (.I(_0267_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1534_ (.A1(_0726_),
    .A2(_0265_),
    .B(_0105_),
    .C(_0778_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1535_ (.A1(_0257_),
    .A2(_0268_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1536_ (.I(_0756_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1537_ (.A1(_0269_),
    .A2(_0680_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1538_ (.I(_0270_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1539_ (.A1(_0709_),
    .A2(_0710_),
    .A3(_0112_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1540_ (.I(_0271_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1541_ (.A1(_0673_),
    .A2(_0254_),
    .B(_0105_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1542_ (.I(_0272_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1543_ (.A1(_0679_),
    .A2(\mod.cpu.state.o_cnt[2] ),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1544_ (.A1(_0679_),
    .A2(\mod.cpu.state.o_cnt[2] ),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1545_ (.A1(_0253_),
    .A2(_0273_),
    .A3(_0274_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1546_ (.A1(_0720_),
    .A2(_0274_),
    .B(_0269_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1547_ (.A1(_0720_),
    .A2(_0274_),
    .B(_0275_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1548_ (.A1(_0720_),
    .A2(_0274_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1549_ (.A1(_0709_),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1550_ (.A1(_0253_),
    .A2(_0277_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1551_ (.A1(_0266_),
    .A2(_0679_),
    .B1(\mod.cpu.i_rf_ready ),
    .B2(_0783_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1552_ (.A1(_0253_),
    .A2(_0278_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1553_ (.A1(_0269_),
    .A2(\mod.cpu.state.o_cnt_r[0] ),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1554_ (.I(_0279_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1555_ (.A1(_0269_),
    .A2(\mod.cpu.state.o_cnt_r[1] ),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1556_ (.I(_0280_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1557_ (.A1(\mod.cpu.mem_bytecnt[1] ),
    .A2(\mod.cpu.bufreg.lsb[1] ),
    .B(\mod.cpu.bufreg.lsb[0] ),
    .C(\mod.cpu.mem_bytecnt[0] ),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1558_ (.A1(\mod.cpu.mem_bytecnt[1] ),
    .A2(\mod.cpu.bufreg.lsb[1] ),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1559_ (.A1(_0603_),
    .A2(_0281_),
    .A3(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1560_ (.A1(_0682_),
    .A2(_0676_),
    .B(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1561_ (.I(_0770_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1562_ (.A1(_0810_),
    .A2(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1563_ (.A1(_0284_),
    .A2(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1564_ (.I(_0285_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1565_ (.A1(_0639_),
    .A2(_0774_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1566_ (.I(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1567_ (.I(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1568_ (.A1(_0812_),
    .A2(_0288_),
    .B(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1569_ (.I(_0776_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1570_ (.A1(_0775_),
    .A2(_0284_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1571_ (.I(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1572_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1573_ (.A1(\mod.cpu.bufreg2.i_dat[0] ),
    .A2(_0293_),
    .B1(_0296_),
    .B2(_0810_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1574_ (.A1(_0287_),
    .A2(_0292_),
    .B(_0297_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1575_ (.I(_0290_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1576_ (.A1(_0814_),
    .A2(_0288_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1577_ (.I(_0284_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1578_ (.A1(\mod.cpu.bufreg2.dat[0] ),
    .A2(_0812_),
    .B(_0285_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1579_ (.A1(_0300_),
    .A2(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1580_ (.I(_0290_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1581_ (.A1(_0812_),
    .A2(_0287_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1582_ (.A1(_0299_),
    .A2(_0302_),
    .B(_0303_),
    .C(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1583_ (.A1(\mod.cpu.bufreg2.i_dat[1] ),
    .A2(_0298_),
    .B(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1584_ (.I(_0306_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1585_ (.A1(\mod.cpu.bufreg2.dat[3] ),
    .A2(_0771_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1586_ (.A1(_0810_),
    .A2(\mod.cpu.bufreg2.dat[1] ),
    .A3(_0814_),
    .B(_0285_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1587_ (.A1(_0300_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1588_ (.A1(_0814_),
    .A2(_0302_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1589_ (.A1(_0307_),
    .A2(_0309_),
    .B(_0303_),
    .C(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1590_ (.A1(\mod.cpu.bufreg2.i_dat[2] ),
    .A2(_0298_),
    .B(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1591_ (.I(_0312_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1592_ (.A1(\mod.cpu.bufreg2.dat[3] ),
    .A2(_0309_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(_0771_),
    .A2(_0767_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1594_ (.A1(_0819_),
    .A2(_0771_),
    .B(_0300_),
    .C(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1595_ (.A1(_0303_),
    .A2(_0313_),
    .A3(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1596_ (.A1(\mod.cpu.bufreg2.i_dat[3] ),
    .A2(_0298_),
    .B(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1597_ (.I(_0317_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1598_ (.A1(_0819_),
    .A2(_0767_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1599_ (.A1(_0288_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1600_ (.A1(_0289_),
    .A2(_0284_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1601_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1602_ (.A1(_0766_),
    .A2(_0288_),
    .B(_0319_),
    .C(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1603_ (.I(_0777_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1604_ (.I(_0294_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1605_ (.I(_0324_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1606_ (.A1(\mod.cpu.bufreg2.i_dat[4] ),
    .A2(_0323_),
    .B1(_0325_),
    .B2(_0819_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1607_ (.A1(_0322_),
    .A2(_0326_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1608_ (.A1(_0290_),
    .A2(_0300_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1609_ (.I(_0295_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1610_ (.A1(\mod.cpu.bufreg2.i_dat[5] ),
    .A2(_0293_),
    .B1(_0328_),
    .B2(_0766_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1611_ (.A1(_0772_),
    .A2(_0327_),
    .B(_0329_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1612_ (.I(_0291_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1613_ (.I(_0324_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1614_ (.I(_0320_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1615_ (.I(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1616_ (.A1(\mod.cpu.bufreg2.dat[6] ),
    .A2(_0331_),
    .B1(_0333_),
    .B2(\mod.cpu.bufreg2.dat[7] ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1617_ (.A1(_1001_),
    .A2(_0330_),
    .B(_0334_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1618_ (.A1(\mod.cpu.bufreg2.dat[7] ),
    .A2(_0331_),
    .B1(_0333_),
    .B2(\mod.cpu.bufreg2.dat[8] ),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1619_ (.A1(_0737_),
    .A2(_0330_),
    .B(_0335_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1620_ (.I(_0776_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1621_ (.I(_0320_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1622_ (.A1(\mod.cpu.bufreg2.i_dat[8] ),
    .A2(_0336_),
    .B1(_0328_),
    .B2(\mod.cpu.bufreg2.dat[8] ),
    .C1(_0337_),
    .C2(\mod.cpu.bufreg2.dat[9] ),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1623_ (.I(_0338_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1624_ (.I(_0777_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1625_ (.A1(\mod.cpu.bufreg2.i_dat[9] ),
    .A2(_0339_),
    .B1(_0328_),
    .B2(\mod.cpu.bufreg2.dat[9] ),
    .C1(_0337_),
    .C2(\mod.cpu.bufreg2.dat[10] ),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1626_ (.I(_0340_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1627_ (.I(_0295_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1628_ (.A1(\mod.cpu.bufreg2.i_dat[10] ),
    .A2(_0339_),
    .B1(_0341_),
    .B2(\mod.cpu.bufreg2.dat[10] ),
    .C1(_0337_),
    .C2(\mod.cpu.bufreg2.dat[11] ),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1629_ (.I(_0342_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1630_ (.A1(\mod.cpu.bufreg2.dat[11] ),
    .A2(_0296_),
    .B1(_0333_),
    .B2(\mod.cpu.bufreg2.dat[12] ),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1631_ (.A1(_0247_),
    .A2(_0330_),
    .B(_0343_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1632_ (.I(_0332_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1633_ (.A1(\mod.cpu.bufreg2.i_dat[12] ),
    .A2(_0339_),
    .B1(_0341_),
    .B2(\mod.cpu.bufreg2.dat[12] ),
    .C1(_0344_),
    .C2(\mod.cpu.bufreg2.dat[13] ),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1634_ (.I(_0345_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1635_ (.A1(\mod.cpu.bufreg2.i_dat[13] ),
    .A2(_0339_),
    .B1(_0341_),
    .B2(\mod.cpu.bufreg2.dat[13] ),
    .C1(_0344_),
    .C2(\mod.cpu.bufreg2.dat[14] ),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1636_ (.I(_0346_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1637_ (.I(_0776_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1638_ (.A1(\mod.cpu.bufreg2.i_dat[14] ),
    .A2(_0347_),
    .B1(_0341_),
    .B2(\mod.cpu.bufreg2.dat[14] ),
    .C1(_0344_),
    .C2(\mod.cpu.bufreg2.dat[15] ),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1639_ (.I(_0348_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1640_ (.I(_0332_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1641_ (.A1(\mod.cpu.bufreg2.dat[16] ),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1642_ (.I(_0324_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1643_ (.A1(\mod.cpu.bufreg2.i_dat[15] ),
    .A2(_0323_),
    .B1(_0351_),
    .B2(\mod.cpu.bufreg2.dat[15] ),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1644_ (.A1(_0350_),
    .A2(_0352_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1645_ (.A1(\mod.cpu.bufreg2.dat[17] ),
    .A2(_0349_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1646_ (.A1(\mod.cpu.bufreg2.i_dat[16] ),
    .A2(_0323_),
    .B1(_0351_),
    .B2(\mod.cpu.bufreg2.dat[16] ),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1647_ (.A1(_0353_),
    .A2(_0354_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1648_ (.I(_0295_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1649_ (.A1(\mod.cpu.bufreg2.i_dat[17] ),
    .A2(_0347_),
    .B1(_0355_),
    .B2(\mod.cpu.bufreg2.dat[17] ),
    .C1(_0344_),
    .C2(\mod.cpu.bufreg2.dat[18] ),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1650_ (.I(_0356_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1651_ (.A1(\mod.cpu.bufreg2.dat[19] ),
    .A2(_0349_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1652_ (.A1(\mod.cpu.bufreg2.i_dat[18] ),
    .A2(_0323_),
    .B1(_0351_),
    .B2(\mod.cpu.bufreg2.dat[18] ),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1653_ (.A1(_0357_),
    .A2(_0358_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1654_ (.I(_0332_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1655_ (.A1(\mod.cpu.bufreg2.i_dat[19] ),
    .A2(_0347_),
    .B1(_0355_),
    .B2(\mod.cpu.bufreg2.dat[19] ),
    .C1(_0359_),
    .C2(\mod.cpu.bufreg2.dat[20] ),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1656_ (.I(_0360_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1657_ (.A1(\mod.cpu.bufreg2.dat[21] ),
    .A2(_0349_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1658_ (.A1(\mod.cpu.bufreg2.i_dat[20] ),
    .A2(_0336_),
    .B1(_0351_),
    .B2(\mod.cpu.bufreg2.dat[20] ),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1659_ (.A1(_0361_),
    .A2(_0362_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1660_ (.A1(\mod.cpu.bufreg2.dat[21] ),
    .A2(_0296_),
    .B1(_0333_),
    .B2(\mod.cpu.bufreg2.dat[22] ),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1661_ (.A1(_0792_),
    .A2(_0330_),
    .B(_0363_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1662_ (.A1(\mod.cpu.bufreg2.i_dat[22] ),
    .A2(_0347_),
    .B1(_0355_),
    .B2(\mod.cpu.bufreg2.dat[22] ),
    .C1(_0359_),
    .C2(\mod.cpu.bufreg2.dat[23] ),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1663_ (.I(_0364_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1664_ (.A1(\mod.cpu.bufreg2.dat[24] ),
    .A2(_0321_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1665_ (.A1(\mod.cpu.bufreg2.i_dat[23] ),
    .A2(_0336_),
    .B1(_0331_),
    .B2(\mod.cpu.bufreg2.dat[23] ),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1666_ (.A1(_0365_),
    .A2(_0366_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1667_ (.A1(\mod.cpu.bufreg2.dat[24] ),
    .A2(_0296_),
    .B1(_0337_),
    .B2(\mod.cpu.bufreg2.dat[25] ),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1668_ (.A1(_0804_),
    .A2(_0298_),
    .B(_0367_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1669_ (.A1(\mod.cpu.bufreg2.i_dat[25] ),
    .A2(_0293_),
    .B1(_0355_),
    .B2(\mod.cpu.bufreg2.dat[25] ),
    .C1(_0359_),
    .C2(\mod.cpu.bufreg2.dat[26] ),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1670_ (.I(_0368_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1671_ (.A1(\mod.cpu.bufreg2.i_dat[26] ),
    .A2(_0291_),
    .B1(_0327_),
    .B2(\mod.cpu.bufreg2.dat[27] ),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1672_ (.A1(_0847_),
    .A2(_0325_),
    .B(_0369_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1673_ (.A1(\mod.cpu.bufreg2.dat[28] ),
    .A2(_0321_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1674_ (.A1(\mod.cpu.bufreg2.i_dat[27] ),
    .A2(_0336_),
    .B1(_0331_),
    .B2(\mod.cpu.bufreg2.dat[27] ),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1675_ (.A1(_0370_),
    .A2(_0371_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1676_ (.A1(\mod.cpu.bufreg2.i_dat[28] ),
    .A2(_0293_),
    .B1(_0324_),
    .B2(\mod.cpu.bufreg2.dat[28] ),
    .C1(_0359_),
    .C2(\mod.cpu.bufreg2.dat[29] ),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1677_ (.I(_0372_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1678_ (.A1(\mod.cpu.bufreg2.i_dat[29] ),
    .A2(_0777_),
    .B1(_0328_),
    .B2(\mod.cpu.bufreg2.dat[29] ),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1679_ (.A1(_0852_),
    .A2(_0327_),
    .B(_0373_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1680_ (.A1(\mod.cpu.bufreg2.i_dat[30] ),
    .A2(_0303_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1681_ (.A1(_0852_),
    .A2(_0325_),
    .B1(_0321_),
    .B2(_0854_),
    .C(_0374_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1682_ (.A1(\mod.cpu.bufreg2.i_dat[31] ),
    .A2(_0291_),
    .B1(_0327_),
    .B2(_0665_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1683_ (.A1(_0854_),
    .A2(_0325_),
    .B(_0375_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1684_ (.A1(_0639_),
    .A2(_0757_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1685_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1686_ (.I(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1687_ (.I(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1688_ (.I(_0376_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1689_ (.A1(\mod.cpu.bufreg2.i_dat[2] ),
    .A2(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1690_ (.A1(_0698_),
    .A2(_0379_),
    .B(_0381_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1691_ (.I(_0376_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1692_ (.I(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1693_ (.I0(_0984_),
    .I1(\mod.cpu.bufreg2.i_dat[3] ),
    .S(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1694_ (.I(_0384_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1695_ (.A1(\mod.cpu.bufreg2.i_dat[4] ),
    .A2(_0380_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1696_ (.A1(_0699_),
    .A2(_0379_),
    .B(_0385_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1697_ (.A1(_0703_),
    .A2(_0759_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1698_ (.A1(_0654_),
    .A2(_0762_),
    .B(_0386_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1699_ (.I(_0759_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1700_ (.I(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1701_ (.A1(_0778_),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1702_ (.A1(_1001_),
    .A2(_0762_),
    .B(_0389_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1703_ (.A1(\mod.cpu.bufreg2.i_dat[12] ),
    .A2(_0382_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1704_ (.A1(_0607_),
    .A2(_0379_),
    .B(_0390_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1705_ (.A1(\mod.cpu.bufreg2.i_dat[13] ),
    .A2(_0382_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1706_ (.A1(_0661_),
    .A2(_0380_),
    .B(_0391_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1707_ (.A1(\mod.cpu.bufreg2.i_dat[14] ),
    .A2(_0382_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1708_ (.I(_0759_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1709_ (.A1(_0658_),
    .A2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1710_ (.A1(_0392_),
    .A2(_0394_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1711_ (.A1(\mod.cpu.bufreg2.i_dat[20] ),
    .A2(_0377_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1712_ (.A1(\mod.cpu.decode.co_ebreak ),
    .A2(_0393_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1713_ (.A1(_0395_),
    .A2(_0396_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1714_ (.I(_0760_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1715_ (.A1(\mod.cpu.immdec.imm24_20[1] ),
    .A2(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1716_ (.A1(_0395_),
    .A2(_0398_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1717_ (.A1(_0726_),
    .A2(_0702_),
    .A3(_0386_),
    .B1(_0376_),
    .B2(_0604_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1718_ (.I0(_0399_),
    .I1(\mod.cpu.immdec.imm24_20[0] ),
    .S(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1719_ (.I(_0401_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1720_ (.I(_0400_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1721_ (.I(_0377_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1722_ (.A1(\mod.cpu.immdec.imm24_20[2] ),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1723_ (.A1(\mod.cpu.bufreg2.i_dat[21] ),
    .A2(_0397_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1724_ (.I(_0400_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1725_ (.A1(\mod.cpu.immdec.imm24_20[1] ),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1726_ (.A1(_0402_),
    .A2(_0404_),
    .A3(_0405_),
    .B(_0407_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1727_ (.A1(\mod.cpu.immdec.imm24_20[3] ),
    .A2(_0387_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1728_ (.A1(\mod.cpu.bufreg2.i_dat[22] ),
    .A2(_0378_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1729_ (.A1(\mod.cpu.immdec.imm24_20[2] ),
    .A2(_0406_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1730_ (.A1(_0402_),
    .A2(_0409_),
    .B(_0410_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1731_ (.A1(\mod.cpu.immdec.imm24_20[4] ),
    .A2(_0387_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1732_ (.A1(\mod.cpu.bufreg2.i_dat[23] ),
    .A2(_0378_),
    .B(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1733_ (.A1(\mod.cpu.immdec.imm24_20[3] ),
    .A2(_0406_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1734_ (.A1(_0402_),
    .A2(_0412_),
    .B(_0413_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1735_ (.A1(\mod.cpu.immdec.imm30_25[0] ),
    .A2(_0387_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1736_ (.A1(\mod.cpu.bufreg2.i_dat[24] ),
    .A2(_0378_),
    .B(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1737_ (.A1(\mod.cpu.immdec.imm24_20[4] ),
    .A2(_0406_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1738_ (.A1(_0402_),
    .A2(_0415_),
    .B(_0416_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1739_ (.A1(_0725_),
    .A2(_0699_),
    .A3(_0704_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1740_ (.A1(_0604_),
    .A2(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1741_ (.I(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1742_ (.I0(\mod.cpu.immdec.imm30_25[1] ),
    .I1(\mod.cpu.immdec.imm30_25[0] ),
    .S(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1743_ (.I(_0758_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1744_ (.I0(\mod.cpu.bufreg2.i_dat[25] ),
    .I1(_0420_),
    .S(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1745_ (.I(_0422_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1746_ (.I0(\mod.cpu.immdec.imm30_25[2] ),
    .I1(\mod.cpu.immdec.imm30_25[1] ),
    .S(_0419_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1747_ (.I(_0760_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1748_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1749_ (.I0(\mod.cpu.bufreg2.i_dat[26] ),
    .I1(_0423_),
    .S(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1750_ (.I(_0426_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1751_ (.I0(\mod.cpu.immdec.imm30_25[3] ),
    .I1(\mod.cpu.immdec.imm30_25[2] ),
    .S(_0418_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1752_ (.I0(\mod.cpu.bufreg2.i_dat[27] ),
    .I1(_0427_),
    .S(_0425_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1753_ (.I(_0428_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1754_ (.I0(\mod.cpu.immdec.imm30_25[4] ),
    .I1(\mod.cpu.immdec.imm30_25[3] ),
    .S(_0418_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1755_ (.I0(\mod.cpu.bufreg2.i_dat[28] ),
    .I1(_0429_),
    .S(_0425_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1756_ (.I(_0430_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1757_ (.I0(\mod.cpu.immdec.imm30_25[5] ),
    .I1(\mod.cpu.immdec.imm30_25[4] ),
    .S(_0418_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1758_ (.I0(\mod.cpu.bufreg2.i_dat[29] ),
    .I1(_0431_),
    .S(_0425_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1759_ (.I(_0432_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1760_ (.I(_0377_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1761_ (.A1(\mod.cpu.bufreg2.i_dat[30] ),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1762_ (.A1(\mod.cpu.immdec.imm31 ),
    .A2(_0620_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1763_ (.A1(_0697_),
    .A2(_0675_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1764_ (.A1(_0984_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1765_ (.I(\mod.cpu.immdec.imm19_12_20[0] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1766_ (.A1(_0438_),
    .A2(_0437_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1767_ (.A1(_0698_),
    .A2(_0729_),
    .B1(_0435_),
    .B2(_0437_),
    .C(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1768_ (.A1(\mod.cpu.immdec.imm7 ),
    .A2(_0986_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1769_ (.A1(_0403_),
    .A2(_0419_),
    .A3(_0440_),
    .A4(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1770_ (.A1(\mod.cpu.immdec.imm30_25[5] ),
    .A2(_0388_),
    .A3(_0419_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1771_ (.A1(_0434_),
    .A2(_0442_),
    .A3(_0443_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1772_ (.A1(\mod.cpu.bufreg2.i_dat[7] ),
    .A2(_0433_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1773_ (.A1(\mod.cpu.immdec.imm7 ),
    .A2(_0783_),
    .A3(_0421_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1774_ (.A1(_0605_),
    .A2(_0435_),
    .A3(_0388_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1775_ (.A1(_0444_),
    .A2(_0445_),
    .A3(_0446_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1776_ (.A1(_0984_),
    .A2(_0682_),
    .B1(_0656_),
    .B2(_0702_),
    .C(_0436_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1777_ (.A1(_0782_),
    .A2(_0447_),
    .B(_0758_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1778_ (.I(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1779_ (.I(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1780_ (.I(_0448_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1781_ (.A1(\mod.cpu.immdec.imm19_12_20[1] ),
    .A2(_0252_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1782_ (.A1(_0395_),
    .A2(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1783_ (.A1(_0451_),
    .A2(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1784_ (.A1(_0438_),
    .A2(_0450_),
    .B(_0454_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1785_ (.A1(\mod.cpu.immdec.imm19_12_20[2] ),
    .A2(_0397_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1786_ (.A1(_0390_),
    .A2(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1787_ (.I(_0448_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1788_ (.I0(\mod.cpu.immdec.imm19_12_20[1] ),
    .I1(_0456_),
    .S(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1789_ (.I(_0458_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1790_ (.A1(\mod.cpu.immdec.imm19_12_20[3] ),
    .A2(_0252_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(_0391_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1792_ (.I0(\mod.cpu.immdec.imm19_12_20[2] ),
    .I1(_0460_),
    .S(_0449_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1793_ (.I(_0461_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1794_ (.A1(\mod.cpu.csr_imm ),
    .A2(_0252_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1795_ (.A1(_0392_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1796_ (.I0(\mod.cpu.immdec.imm19_12_20[3] ),
    .I1(_0463_),
    .S(_0449_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1797_ (.I(_0464_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1798_ (.A1(\mod.cpu.immdec.imm19_12_20[5] ),
    .A2(_0424_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1799_ (.A1(\mod.cpu.bufreg2.i_dat[15] ),
    .A2(_0383_),
    .B(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1800_ (.A1(\mod.cpu.csr_imm ),
    .A2(_0451_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1801_ (.A1(_0450_),
    .A2(_0466_),
    .B(_0467_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1802_ (.A1(\mod.cpu.immdec.imm19_12_20[6] ),
    .A2(_0424_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1803_ (.A1(\mod.cpu.bufreg2.i_dat[16] ),
    .A2(_0383_),
    .B(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1804_ (.A1(\mod.cpu.immdec.imm19_12_20[5] ),
    .A2(_0457_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1805_ (.A1(_0450_),
    .A2(_0469_),
    .B(_0470_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1806_ (.A1(\mod.cpu.immdec.imm19_12_20[7] ),
    .A2(_0424_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1807_ (.A1(\mod.cpu.bufreg2.i_dat[17] ),
    .A2(_0433_),
    .B(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1808_ (.A1(\mod.cpu.immdec.imm19_12_20[6] ),
    .A2(_0457_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1809_ (.A1(_0451_),
    .A2(_0472_),
    .B(_0473_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1810_ (.A1(_0645_),
    .A2(_0403_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1811_ (.A1(\mod.cpu.bufreg2.i_dat[18] ),
    .A2(_0433_),
    .B(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1812_ (.A1(\mod.cpu.immdec.imm19_12_20[7] ),
    .A2(_0457_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1813_ (.A1(_0451_),
    .A2(_0475_),
    .B(_0476_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1814_ (.A1(_0701_),
    .A2(\mod.cpu.immdec.imm24_20[0] ),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1815_ (.A1(_0778_),
    .A2(_0435_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1816_ (.A1(_0397_),
    .A2(_0477_),
    .A3(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1817_ (.A1(\mod.cpu.bufreg2.i_dat[19] ),
    .A2(_0421_),
    .B(_0449_),
    .C(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1818_ (.A1(_0645_),
    .A2(_0450_),
    .B(_0480_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1819_ (.I0(\mod.cpu.immdec.imm31 ),
    .I1(\mod.cpu.bufreg2.i_dat[31] ),
    .S(_0383_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1820_ (.I(_0481_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1821_ (.A1(\mod.cpu.bufreg.i_sh_signed ),
    .A2(_0388_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1822_ (.A1(_0434_),
    .A2(_0482_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1823_ (.I0(\mod.cpu.alu.cmp_r ),
    .I1(_0264_),
    .S(_0605_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1824_ (.I(_0483_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1825_ (.I(_0692_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1826_ (.I(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1827_ (.I0(\mod.cpu.bufreg.data[2] ),
    .I1(\mod.cpu.bufreg.data[3] ),
    .S(_0485_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1828_ (.I(_0486_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1829_ (.I0(\mod.cpu.bufreg.data[3] ),
    .I1(\mod.cpu.bufreg.data[4] ),
    .S(_0485_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1830_ (.I(_0487_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1831_ (.I0(\mod.cpu.bufreg.data[4] ),
    .I1(\mod.cpu.bufreg.data[5] ),
    .S(_0485_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1832_ (.I(_0488_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1833_ (.I0(\mod.cpu.bufreg.data[5] ),
    .I1(\mod.cpu.bufreg.data[6] ),
    .S(_0485_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1834_ (.I(_0489_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1835_ (.I(_0484_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1836_ (.I0(\mod.cpu.bufreg.data[6] ),
    .I1(\mod.cpu.bufreg.data[7] ),
    .S(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1837_ (.I(_0491_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1838_ (.I0(\mod.cpu.bufreg.data[7] ),
    .I1(\mod.cpu.bufreg.data[8] ),
    .S(_0490_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1839_ (.I(_0492_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1840_ (.I0(\mod.cpu.bufreg.data[8] ),
    .I1(\mod.cpu.bufreg.data[9] ),
    .S(_0490_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1841_ (.I(_0493_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1842_ (.I0(\mod.cpu.bufreg.data[9] ),
    .I1(\mod.cpu.bufreg.data[10] ),
    .S(_0490_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1843_ (.I(_0494_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1844_ (.I(_0692_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1845_ (.I(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1846_ (.I0(\mod.cpu.bufreg.data[10] ),
    .I1(\mod.cpu.bufreg.data[11] ),
    .S(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1847_ (.I(_0497_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1848_ (.I0(\mod.cpu.bufreg.data[11] ),
    .I1(\mod.cpu.bufreg.data[12] ),
    .S(_0496_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1849_ (.I(_0498_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1850_ (.I0(\mod.cpu.bufreg.data[12] ),
    .I1(\mod.cpu.bufreg.data[13] ),
    .S(_0496_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1851_ (.I(_0499_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1852_ (.I0(\mod.cpu.bufreg.data[13] ),
    .I1(\mod.cpu.bufreg.data[14] ),
    .S(_0496_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1853_ (.I(_0500_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1854_ (.I(_0495_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1855_ (.I0(\mod.cpu.bufreg.data[14] ),
    .I1(\mod.cpu.bufreg.data[15] ),
    .S(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1856_ (.I(_0502_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1857_ (.I0(\mod.cpu.bufreg.data[15] ),
    .I1(\mod.cpu.bufreg.data[16] ),
    .S(_0501_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1858_ (.I(_0503_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1859_ (.I0(\mod.cpu.bufreg.data[16] ),
    .I1(\mod.cpu.bufreg.data[17] ),
    .S(_0501_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1860_ (.I(_0504_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1861_ (.I0(\mod.cpu.bufreg.data[17] ),
    .I1(\mod.cpu.bufreg.data[18] ),
    .S(_0501_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1862_ (.I(_0505_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1863_ (.I(_0495_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1864_ (.I0(\mod.cpu.bufreg.data[18] ),
    .I1(\mod.cpu.bufreg.data[19] ),
    .S(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1865_ (.I(_0507_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1866_ (.I0(\mod.cpu.bufreg.data[19] ),
    .I1(\mod.cpu.bufreg.data[20] ),
    .S(_0506_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1867_ (.I(_0508_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1868_ (.I0(\mod.cpu.bufreg.data[20] ),
    .I1(\mod.cpu.bufreg.data[21] ),
    .S(_0506_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1869_ (.I(_0509_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1870_ (.I0(\mod.cpu.bufreg.data[21] ),
    .I1(\mod.cpu.bufreg.data[22] ),
    .S(_0506_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1871_ (.I(_0510_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1872_ (.I(_0495_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1873_ (.I0(\mod.cpu.bufreg.data[22] ),
    .I1(\mod.cpu.bufreg.data[23] ),
    .S(_0511_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1874_ (.I(_0512_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1875_ (.I0(\mod.cpu.bufreg.data[23] ),
    .I1(\mod.cpu.bufreg.data[24] ),
    .S(_0511_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1876_ (.I(_0513_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1877_ (.I0(\mod.cpu.bufreg.data[24] ),
    .I1(\mod.cpu.bufreg.data[25] ),
    .S(_0511_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1878_ (.I(_0514_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1879_ (.I0(\mod.cpu.bufreg.data[25] ),
    .I1(\mod.cpu.bufreg.data[26] ),
    .S(_0511_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1880_ (.I(_0515_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1881_ (.I(_0692_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1882_ (.I0(\mod.cpu.bufreg.data[26] ),
    .I1(\mod.cpu.bufreg.data[27] ),
    .S(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1883_ (.I(_0517_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1884_ (.I0(\mod.cpu.bufreg.data[27] ),
    .I1(\mod.cpu.bufreg.data[28] ),
    .S(_0516_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1885_ (.I(_0518_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1886_ (.I0(\mod.cpu.bufreg.data[28] ),
    .I1(\mod.cpu.bufreg.data[29] ),
    .S(_0516_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1887_ (.I(_0519_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1888_ (.I0(\mod.cpu.bufreg.data[29] ),
    .I1(\mod.cpu.bufreg.data[30] ),
    .S(_0516_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1889_ (.I(_0520_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1890_ (.I0(\mod.cpu.bufreg.data[30] ),
    .I1(\mod.cpu.bufreg.data[31] ),
    .S(_0484_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1891_ (.I(_0521_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1892_ (.I(_0764_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1893_ (.A1(_0989_),
    .A2(_0992_),
    .B(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1894_ (.A1(_0989_),
    .A2(_0992_),
    .B(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1895_ (.A1(\mod.cpu.bufreg.i_sh_signed ),
    .A2(\mod.cpu.bufreg.data[31] ),
    .A3(_0522_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1896_ (.A1(_0524_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1897_ (.I0(\mod.cpu.bufreg.data[31] ),
    .I1(_0526_),
    .S(_0484_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1898_ (.I(_0527_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1899_ (.A1(_0602_),
    .A2(_0730_),
    .B(_0764_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1900_ (.A1(_0522_),
    .A2(_0996_),
    .B(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1901_ (.A1(_0806_),
    .A2(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1902_ (.A1(_0805_),
    .A2(_0529_),
    .B(_0530_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1903_ (.A1(\mod.cpu.bufreg.data[2] ),
    .A2(_0522_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1904_ (.A1(_0524_),
    .A2(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1905_ (.I0(_0806_),
    .I1(_0532_),
    .S(_0529_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1906_ (.I(_0533_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1907_ (.A1(_0249_),
    .A2(_0740_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1908_ (.I(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1909_ (.I(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1910_ (.A1(_0859_),
    .A2(_0251_),
    .B1(_0536_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[1] ),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1911_ (.I(_0537_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1912_ (.A1(\mod.cpu.ctrl.o_ibus_adr[1] ),
    .A2(_0251_),
    .B1(_0536_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1913_ (.I(_0538_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1914_ (.I(_0250_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1915_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1916_ (.A1(\mod.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_0540_),
    .B1(_0536_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1917_ (.I(_0541_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1918_ (.A1(\mod.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0540_),
    .B1(_0536_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1919_ (.I(_0542_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1920_ (.I(_0535_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1921_ (.A1(\mod.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0540_),
    .B1(_0543_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[5] ),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1922_ (.I(_0544_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1923_ (.A1(\mod.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_0540_),
    .B1(_0543_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1924_ (.I(_0545_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1925_ (.I(_0539_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1926_ (.A1(\mod.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_0546_),
    .B1(_0543_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1927_ (.I(_0547_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1928_ (.A1(\mod.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0546_),
    .B1(_0543_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1929_ (.I(_0548_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1930_ (.I(_0535_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1931_ (.A1(\mod.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_0546_),
    .B1(_0549_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1932_ (.I(_0550_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1933_ (.A1(\mod.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0546_),
    .B1(_0549_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1934_ (.I(_0551_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1935_ (.I(_0539_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1936_ (.A1(\mod.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0552_),
    .B1(_0549_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1937_ (.I(_0553_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1938_ (.A1(\mod.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_0552_),
    .B1(_0549_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[12] ),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1939_ (.I(_0554_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1940_ (.I(_0535_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1941_ (.A1(\mod.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_0552_),
    .B1(_0555_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1942_ (.I(_0556_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1943_ (.A1(\mod.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_0552_),
    .B1(_0555_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1944_ (.I(_0557_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1945_ (.I(_0250_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1946_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1947_ (.A1(\mod.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0559_),
    .B1(_0555_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1948_ (.I(_0560_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1949_ (.A1(\mod.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_0559_),
    .B1(_0555_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1950_ (.I(_0561_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1951_ (.I(_0534_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1952_ (.I(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1953_ (.A1(\mod.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0559_),
    .B1(_0563_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1954_ (.I(_0564_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1955_ (.A1(\mod.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_0559_),
    .B1(_0563_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1956_ (.I(_0565_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1957_ (.I(_0558_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1958_ (.A1(\mod.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0566_),
    .B1(_0563_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1959_ (.I(_0567_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1960_ (.A1(\mod.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_0566_),
    .B1(_0563_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1961_ (.I(_0568_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1962_ (.I(_0562_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1963_ (.A1(\mod.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0566_),
    .B1(_0569_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1964_ (.I(_0570_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1965_ (.A1(\mod.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0566_),
    .B1(_0569_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1966_ (.I(_0571_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1967_ (.I(_0558_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1968_ (.A1(\mod.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0572_),
    .B1(_0569_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1969_ (.I(_0573_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1970_ (.A1(\mod.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0572_),
    .B1(_0569_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1971_ (.I(_0574_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1972_ (.I(_0562_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1973_ (.A1(\mod.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_0572_),
    .B1(_0575_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1974_ (.I(_0576_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1975_ (.A1(\mod.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0572_),
    .B1(_0575_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1976_ (.I(_0577_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1977_ (.I(_0558_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1978_ (.A1(\mod.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0578_),
    .B1(_0575_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1979_ (.I(_0579_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1980_ (.A1(\mod.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_0578_),
    .B1(_0575_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1981_ (.I(_0580_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1982_ (.I(_0562_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1983_ (.A1(\mod.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0578_),
    .B1(_0581_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1984_ (.I(_0582_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1985_ (.A1(\mod.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0578_),
    .B1(_0581_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1986_ (.I(_0583_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1987_ (.A1(\mod.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_0539_),
    .B1(_0581_),
    .B2(\mod.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1988_ (.I(_0584_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1989_ (.A1(\mod.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0251_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1990_ (.A1(\mod.cpu.ctrl.i_jump ),
    .A2(_0716_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1991_ (.A1(\mod.cpu.ctrl.i_jump ),
    .A2(_0733_),
    .B(_0581_),
    .C(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1992_ (.A1(_0585_),
    .A2(_0587_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1993_ (.A1(_0782_),
    .A2(_0743_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1994_ (.I0(\mod.cpu.immdec.imm11_7[0] ),
    .I1(\mod.cpu.immdec.imm11_7[1] ),
    .S(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1995_ (.A1(_0393_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1996_ (.A1(_0444_),
    .A2(_0590_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1997_ (.I(_0588_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1998_ (.I(_0588_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1999_ (.A1(_0747_),
    .A2(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2000_ (.A1(\mod.cpu.immdec.imm11_7[1] ),
    .A2(_0591_),
    .B(_0593_),
    .C(_0761_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2001_ (.A1(_1003_),
    .A2(_0762_),
    .B(_0594_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2002_ (.A1(_0751_),
    .A2(_0592_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2003_ (.A1(\mod.cpu.immdec.imm11_7[2] ),
    .A2(_0591_),
    .B(_0595_),
    .C(_0761_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2004_ (.A1(_1004_),
    .A2(_0393_),
    .B(_0596_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2005_ (.A1(_0751_),
    .A2(_0592_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2006_ (.A1(\mod.cpu.immdec.imm11_7[4] ),
    .A2(_0592_),
    .B(_0597_),
    .C(_0403_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2007_ (.A1(_1005_),
    .A2(_0379_),
    .B(_0598_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2008_ (.A1(\mod.cpu.immdec.imm11_7[4] ),
    .A2(_0761_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2009_ (.A1(\mod.cpu.bufreg2.i_dat[11] ),
    .A2(_0380_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2010_ (.A1(\mod.cpu.immdec.imm30_25[0] ),
    .A2(_0421_),
    .A3(_0591_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2011_ (.A1(_0591_),
    .A2(_0599_),
    .B(_0600_),
    .C(_0601_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2012_ (.D(_0004_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_rs2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2013_ (.D(_0008_),
    .CLK(net4),
    .Q(\mod.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2014_ (.D(_0019_),
    .CLK(net4),
    .Q(\mod.cpu.i_rf_ready ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2015_ (.D(_0030_),
    .CLK(net4),
    .Q(\mod.cpu.i_timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2016_ (.D(_0041_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2017_ (.D(_0052_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2018_ (.D(_0063_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2019_ (.D(_0074_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2020_ (.D(_0085_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2021_ (.D(_0092_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2022_ (.D(_0005_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2023_ (.D(_0006_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2024_ (.D(_0007_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2025_ (.D(_0009_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2026_ (.D(_0010_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2027_ (.D(_0011_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2028_ (.D(_0012_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2029_ (.D(_0013_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2030_ (.D(_0014_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2031_ (.D(_0015_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2032_ (.D(_0016_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2033_ (.D(_0017_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2034_ (.D(_0018_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2035_ (.D(_0020_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2036_ (.D(_0021_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2037_ (.D(_0022_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2038_ (.D(_0023_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2039_ (.D(_0024_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2040_ (.D(_0025_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2041_ (.D(_0026_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2042_ (.D(_0027_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2043_ (.D(_0028_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2044_ (.D(_0029_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2045_ (.D(_0031_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2046_ (.D(_0032_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2047_ (.D(_0033_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2048_ (.D(_0034_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2049_ (.D(_0035_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2050_ (.D(_0036_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2051_ (.D(_0037_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2052_ (.D(_0038_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2053_ (.D(_0039_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2054_ (.D(_0040_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2055_ (.D(_0042_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2056_ (.D(_0043_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2057_ (.D(_0044_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2058_ (.D(_0045_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2059_ (.D(_0046_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2060_ (.D(_0047_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2061_ (.D(_0048_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2062_ (.D(_0049_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2063_ (.D(_0050_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2064_ (.D(_0051_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2065_ (.D(_0053_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2066_ (.D(_0054_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2067_ (.D(_0055_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2068_ (.D(_0056_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2069_ (.D(_0057_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2070_ (.D(_0058_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2071_ (.D(_0059_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2072_ (.D(_0060_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2073_ (.D(_0061_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2074_ (.D(_0062_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2075_ (.D(_0064_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2076_ (.D(_0065_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2077_ (.D(_0066_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2078_ (.D(_0067_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2079_ (.D(_0068_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2080_ (.D(_0069_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2081_ (.D(_0070_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2082_ (.D(_0071_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2083_ (.D(_0072_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2084_ (.D(_0073_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2085_ (.D(_0075_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[80] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2086_ (.D(_0076_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[81] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2087_ (.D(_0077_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[82] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2088_ (.D(_0078_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[83] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2089_ (.D(_0079_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[84] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2090_ (.D(_0080_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[85] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2091_ (.D(_0081_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[86] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2092_ (.D(_0082_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[87] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2093_ (.D(_0083_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[88] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2094_ (.D(_0084_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[89] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2095_ (.D(_0086_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[90] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2096_ (.D(_0087_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[91] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2097_ (.D(_0088_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[92] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2098_ (.D(_0089_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[93] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2099_ (.D(_0090_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[94] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2100_ (.D(_0091_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[95] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2101_ (.D(_0093_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2102_ (.D(_0094_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2103_ (.D(_0095_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2104_ (.D(_0096_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2105_ (.D(_0097_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2106_ (.D(_0098_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2107_ (.D(_0099_),
    .CLK(net4),
    .Q(\mod.cpu.bufreg2.i_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2108_ (.D(_0100_),
    .CLK(net3),
    .Q(\mod.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _2109_ (.D(\mod.u_scanchain_local.module_data_in[95] ),
    .CLKN(net4),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2110_ (.D(_0101_),
    .CLK(net3),
    .Q(\mod.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2111_ (.D(_0102_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2112_ (.D(_0103_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2113_ (.D(_0104_),
    .CLK(net3),
    .Q(\mod.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2114_ (.D(_0105_),
    .CLK(net3),
    .Q(\mod.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2115_ (.D(_0106_),
    .CLK(net3),
    .Q(\mod.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2116_ (.D(_0107_),
    .CLK(net3),
    .Q(\mod.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2117_ (.D(_0108_),
    .CLK(net3),
    .Q(\mod.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2118_ (.D(_0109_),
    .CLK(net3),
    .Q(\mod.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2119_ (.D(_0110_),
    .CLK(net3),
    .Q(\mod.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2120_ (.D(_0111_),
    .CLK(net3),
    .Q(\mod.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2121_ (.D(_0112_),
    .CLK(net3),
    .Q(\mod.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2122_ (.D(_0113_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2123_ (.D(_0114_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2124_ (.D(_0115_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2125_ (.D(_0116_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2126_ (.D(_0117_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2127_ (.D(_0118_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2128_ (.D(_0119_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2129_ (.D(_0120_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2130_ (.D(_0121_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2131_ (.D(_0122_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2132_ (.D(_0123_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2133_ (.D(_0124_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2134_ (.D(_0125_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2135_ (.D(_0126_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2136_ (.D(_0127_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2137_ (.D(_0128_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2138_ (.D(_0129_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2139_ (.D(_0130_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2140_ (.D(_0131_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2141_ (.D(_0132_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2142_ (.D(_0133_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2143_ (.D(_0134_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2144_ (.D(_0135_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2145_ (.D(_0136_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2146_ (.D(_0137_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2147_ (.D(_0138_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2148_ (.D(_0139_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2149_ (.D(_0140_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2150_ (.D(_0141_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2151_ (.D(_0142_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2152_ (.D(_0143_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2153_ (.D(_0144_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2154_ (.D(_0145_),
    .CLK(net3),
    .Q(\mod.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2155_ (.D(_0146_),
    .CLK(net3),
    .Q(\mod.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2156_ (.D(_0147_),
    .CLK(net3),
    .Q(\mod.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2157_ (.D(_0148_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg2.i_op_b_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2158_ (.D(_0149_),
    .CLK(net3),
    .Q(\mod.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2159_ (.D(_0150_),
    .CLK(net3),
    .Q(\mod.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2160_ (.D(_0151_),
    .CLK(net3),
    .Q(\mod.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2161_ (.D(_0152_),
    .CLK(net3),
    .Q(\mod.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2162_ (.D(_0153_),
    .CLK(net3),
    .Q(\mod.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2163_ (.D(_0154_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2164_ (.D(_0155_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2165_ (.D(_0156_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2166_ (.D(_0157_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2167_ (.D(_0158_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2168_ (.D(_0159_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2169_ (.D(_0160_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2170_ (.D(_0161_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2171_ (.D(_0162_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2172_ (.D(_0163_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2173_ (.D(_0164_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2174_ (.D(_0165_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2175_ (.D(_0166_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2176_ (.D(_0167_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2177_ (.D(_0168_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2178_ (.D(_0169_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2179_ (.D(_0170_),
    .CLK(net3),
    .Q(\mod.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2180_ (.D(_0171_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2181_ (.D(_0172_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2182_ (.D(_0173_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2183_ (.D(_0174_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2184_ (.D(_0175_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2185_ (.D(_0176_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2186_ (.D(_0177_),
    .CLK(net3),
    .Q(\mod.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2187_ (.D(_0178_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2188_ (.D(_0179_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2189_ (.D(_0180_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2190_ (.D(_0181_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2191_ (.D(_0182_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2192_ (.D(_0183_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2193_ (.D(_0184_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2194_ (.D(_0185_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2195_ (.D(_0186_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2196_ (.D(_0187_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2197_ (.D(_0188_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2198_ (.D(_0189_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2199_ (.D(_0190_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2200_ (.D(_0191_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2201_ (.D(_0192_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2202_ (.D(_0193_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2203_ (.D(_0194_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2204_ (.D(_0195_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2205_ (.D(_0196_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2206_ (.D(_0197_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2207_ (.D(_0198_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2208_ (.D(_0199_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2209_ (.D(_0200_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2210_ (.D(_0201_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2211_ (.D(_0202_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2212_ (.D(_0203_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2213_ (.D(_0204_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2214_ (.D(_0205_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2215_ (.D(_0206_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2216_ (.D(_0207_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2217_ (.D(_0001_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2218_ (.D(_0208_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2219_ (.D(_0209_),
    .CLK(net3),
    .Q(\mod.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2220_ (.D(_0003_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2221_ (.D(_0002_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2222_ (.D(_0210_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2223_ (.D(_0211_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2224_ (.D(_0212_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2225_ (.D(_0213_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2226_ (.D(_0214_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2227_ (.D(_0215_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2228_ (.D(_0216_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2229_ (.D(_0217_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2230_ (.D(_0218_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2231_ (.D(_0219_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2232_ (.D(_0220_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2233_ (.D(_0221_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2234_ (.D(_0222_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2235_ (.D(_0223_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2236_ (.D(_0224_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2237_ (.D(_0225_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2238_ (.D(_0226_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2239_ (.D(_0227_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2240_ (.D(_0228_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2241_ (.D(_0229_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2242_ (.D(_0230_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2243_ (.D(_0231_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2244_ (.D(_0232_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2245_ (.D(_0233_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2246_ (.D(_0234_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2247_ (.D(_0235_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2248_ (.D(_0236_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2249_ (.D(_0237_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2250_ (.D(_0238_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2251_ (.D(_0239_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2252_ (.D(_0240_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2253_ (.D(_0241_),
    .CLK(net3),
    .Q(\mod.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2254_ (.D(_0000_),
    .CLK(net3),
    .Q(\mod.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2255_ (.D(_0242_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2256_ (.D(_0243_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2257_ (.D(_0244_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2258_ (.D(_0245_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2259_ (.D(_0246_),
    .CLK(net3),
    .Q(\mod.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_9 (.ZN(net9));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_10 (.ZN(net10));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_11 (.ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_12 (.ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_13 (.ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_14 (.ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_15 (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__D (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2433_ (.I(net4),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2434_ (.I(net2),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[12]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[13]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input3 (.I(io_in[15]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 input4 (.I(io_in[8]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output5 (.I(net5),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output6 (.I(net6),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output7 (.I(net7),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_8 (.ZN(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__D (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A2 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__A2 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A2 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__B (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__I (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__B (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__B (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__I (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__I (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__B (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__B1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__B (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__B (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__B1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__C (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__B1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__I (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__I (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__I (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__B1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__B1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__B1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__B1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__B1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__B1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__B1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__B1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__B1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__B1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__B1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__C1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__C1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__C1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__C1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__C1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__C1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__C1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__B1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__S (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__S (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A3 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__B (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__I (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__I (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__S (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__C (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__S (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__S (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__S (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A3 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__S (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__S (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A3 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__S (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__S (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__S (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__S (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__S (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__B (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__S (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__S (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__I (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__S (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__S (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__S (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__I (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__I (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__S (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__S (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__S (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__S (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__S (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__S (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__S (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__S (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__I1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__B (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__B1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__B1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__B1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__B2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__S (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1033__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1136__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1026__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1104__B (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1070__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1126__B (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1027__I1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1250__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1144__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1035__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1215__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1046__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1042__I0 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__S (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__S (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__S (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1047__S (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1199__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__I0 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1068__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1435__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1062__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1168__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1320__I (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1169__I (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__I (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1318__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1314__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1153__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__B1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1087__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1072__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1197__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1197__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1079__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1486__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1131__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1079__A3 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__B2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1085__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1083__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__A3 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1084__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1093__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1114__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1092__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1096__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1128__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1109__C (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1115__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1152__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1128__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1127__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1486__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1160__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1119__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A3 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1122__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1140__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1140__A3 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1225__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__S1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1150__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__B (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1225__B (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1161__C (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1151__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1150__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1496__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1147__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1150__A3 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1194__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1188__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__B (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__B (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__B1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1161__B (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1171__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1173__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1427__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1317__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1323__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1181__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1183__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__B (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__I (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A3 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1196__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1197__A3 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1199__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1203__B (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__C (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1203__C (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__I (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__S (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__S (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__B2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__A3 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__A3 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1210__B (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1410__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1214__B (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__I1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__S (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__S (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__S (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__S (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1328__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1231__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__A3 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__B (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A3 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__I1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1279__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1270__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1261__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1251__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__S (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__S (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__S (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__S (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1286__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1284__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__S (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1293__S (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__S (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1289__S (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__S (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1302__S (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1300__S (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1298__S (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1344__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1319__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1327__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1341__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1324__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1333__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__B (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__B (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__B (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__B (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1411__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1436__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__I0 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A3 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A4 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1102__A2 (.I(\mod.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__I (.I(\mod.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A2 (.I(\mod.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__C (.I(\mod.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__I0 (.I(\mod.cpu.bufreg.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__I1 (.I(\mod.cpu.bufreg.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A1 (.I(\mod.cpu.bufreg.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__I0 (.I(\mod.cpu.bufreg.data[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I1 (.I(\mod.cpu.bufreg.data[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A1 (.I(\mod.cpu.bufreg.data[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A1 (.I(\mod.cpu.bufreg.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__I0 (.I(\mod.cpu.bufreg.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__A1 (.I(\mod.cpu.bufreg.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__I0 (.I(\mod.cpu.bufreg.data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A2 (.I(\mod.cpu.bufreg.data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__I1 (.I(\mod.cpu.bufreg.data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A1 (.I(\mod.cpu.bufreg.data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__I0 (.I(\mod.cpu.bufreg.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__I1 (.I(\mod.cpu.bufreg.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A1 (.I(\mod.cpu.bufreg.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(\mod.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A1 (.I(\mod.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__A2 (.I(\mod.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__B (.I(\mod.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1224__I (.I(\mod.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__S0 (.I(\mod.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__A1 (.I(\mod.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A2 (.I(\mod.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__A2 (.I(\mod.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__I (.I(\mod.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A1 (.I(\mod.cpu.bufreg2.dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__I (.I(\mod.cpu.bufreg2.dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__A1 (.I(\mod.cpu.bufreg2.dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__I0 (.I(\mod.cpu.bufreg2.dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__B2 (.I(\mod.cpu.bufreg2.dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__C2 (.I(\mod.cpu.bufreg2.dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__I1 (.I(\mod.cpu.bufreg2.dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A1 (.I(\mod.cpu.bufreg2.dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__C2 (.I(\mod.cpu.bufreg2.dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1271__I1 (.I(\mod.cpu.bufreg2.dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__B2 (.I(\mod.cpu.bufreg2.dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__B2 (.I(\mod.cpu.bufreg2.dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__I1 (.I(\mod.cpu.bufreg2.dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__B2 (.I(\mod.cpu.bufreg2.dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__C2 (.I(\mod.cpu.bufreg2.dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1277__I1 (.I(\mod.cpu.bufreg2.dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__B2 (.I(\mod.cpu.bufreg2.dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(\mod.cpu.bufreg2.dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__I1 (.I(\mod.cpu.bufreg2.dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__I2 (.I(\mod.cpu.bufreg2.dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B2 (.I(\mod.cpu.bufreg2.dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A1 (.I(\mod.cpu.bufreg2.dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1289__I1 (.I(\mod.cpu.bufreg2.dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A1 (.I(\mod.cpu.bufreg2.dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A1 (.I(\mod.cpu.bufreg2.dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1293__I1 (.I(\mod.cpu.bufreg2.dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__B2 (.I(\mod.cpu.bufreg2.dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__B2 (.I(\mod.cpu.bufreg2.dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__I1 (.I(\mod.cpu.bufreg2.dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__B2 (.I(\mod.cpu.bufreg2.dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__C2 (.I(\mod.cpu.bufreg2.dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1298__I1 (.I(\mod.cpu.bufreg2.dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(\mod.cpu.bufreg2.dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A1 (.I(\mod.cpu.bufreg2.dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1300__I1 (.I(\mod.cpu.bufreg2.dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__I3 (.I(\mod.cpu.bufreg2.dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__B2 (.I(\mod.cpu.bufreg2.dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B2 (.I(\mod.cpu.bufreg2.dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1302__I1 (.I(\mod.cpu.bufreg2.dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__B2 (.I(\mod.cpu.bufreg2.dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__B2 (.I(\mod.cpu.bufreg2.dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__I1 (.I(\mod.cpu.bufreg2.dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__B2 (.I(\mod.cpu.bufreg2.dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A1 (.I(\mod.cpu.bufreg2.dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__I1 (.I(\mod.cpu.bufreg2.dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__B2 (.I(\mod.cpu.bufreg2.dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__C2 (.I(\mod.cpu.bufreg2.dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__I1 (.I(\mod.cpu.bufreg2.dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1190__I (.I(\mod.cpu.bufreg2.dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1087__A2 (.I(\mod.cpu.bufreg2.dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(\mod.cpu.bufreg2.dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__I1 (.I(\mod.cpu.bufreg2.dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1196__A1 (.I(\mod.cpu.bufreg2.dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A1 (.I(\mod.cpu.bufreg2.dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__B2 (.I(\mod.cpu.bufreg2.dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__I1 (.I(\mod.cpu.bufreg2.dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__B2 (.I(\mod.cpu.bufreg2.dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__B2 (.I(\mod.cpu.bufreg2.dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__I1 (.I(\mod.cpu.bufreg2.dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__I1 (.I(\mod.cpu.bufreg2.dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__B2 (.I(\mod.cpu.bufreg2.dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__C2 (.I(\mod.cpu.bufreg2.dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__I1 (.I(\mod.cpu.bufreg2.dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__A1 (.I(\mod.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1016__I (.I(\mod.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A1 (.I(\mod.cpu.bufreg2.i_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__I0 (.I(\mod.cpu.bufreg2.i_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(\mod.cpu.bufreg2.i_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__I (.I(\mod.cpu.bufreg2.i_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A1 (.I(\mod.cpu.bufreg2.i_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__I (.I(\mod.cpu.bufreg2.i_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A1 (.I(\mod.cpu.bufreg2.i_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A1 (.I(\mod.cpu.bufreg2.i_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A1 (.I(\mod.cpu.bufreg2.i_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A1 (.I(\mod.cpu.bufreg2.i_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__A1 (.I(\mod.cpu.bufreg2.i_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__I0 (.I(\mod.cpu.bufreg2.i_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(\mod.cpu.bufreg2.i_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A1 (.I(\mod.cpu.bufreg2.i_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__I0 (.I(\mod.cpu.bufreg2.i_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A1 (.I(\mod.cpu.bufreg2.i_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A1 (.I(\mod.cpu.bufreg2.i_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__A1 (.I(\mod.cpu.bufreg2.i_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A1 (.I(\mod.cpu.bufreg2.i_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A1 (.I(\mod.cpu.bufreg2.i_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1173__A1 (.I(\mod.cpu.bufreg2.i_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A1 (.I(\mod.cpu.bufreg2.i_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(\mod.cpu.bufreg2.i_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__I0 (.I(\mod.cpu.bufreg2.i_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(\mod.cpu.bufreg2.i_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A1 (.I(\mod.cpu.bufreg2.i_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__A1 (.I(\mod.cpu.bufreg2.i_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A1 (.I(\mod.cpu.bufreg2.i_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(\mod.cpu.bufreg2.i_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__A1 (.I(\mod.cpu.bufreg2.i_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(\mod.cpu.bufreg2.i_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__I0 (.I(\mod.cpu.bufreg2.i_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(\mod.cpu.bufreg2.i_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(\mod.cpu.bufreg2.i_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__I0 (.I(\mod.cpu.bufreg2.i_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(\mod.cpu.bufreg2.i_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1218__I (.I(\mod.cpu.bufreg2.i_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(\mod.cpu.bufreg2.i_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A1 (.I(\mod.cpu.bufreg2.i_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__A1 (.I(\mod.cpu.bufreg2.i_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A1 (.I(\mod.cpu.bufreg2.i_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A1 (.I(\mod.cpu.bufreg2.i_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1231__A1 (.I(\mod.cpu.bufreg2.i_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A1 (.I(\mod.cpu.bufreg2.i_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1233__I (.I(\mod.cpu.bufreg2.i_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__I0 (.I(\mod.cpu.bufreg2.i_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(\mod.cpu.bufreg2.i_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__I (.I(\mod.cpu.bufreg2.i_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__I0 (.I(\mod.cpu.bufreg2.i_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__A1 (.I(\mod.cpu.bufreg2.i_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__I0 (.I(\mod.cpu.bufreg2.i_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__I0 (.I(\mod.cpu.bufreg2.i_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A1 (.I(\mod.cpu.bufreg2.i_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__I0 (.I(\mod.cpu.bufreg2.i_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__I0 (.I(\mod.cpu.bufreg2.i_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A1 (.I(\mod.cpu.bufreg2.i_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__I0 (.I(\mod.cpu.bufreg2.i_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__I0 (.I(\mod.cpu.bufreg2.i_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A1 (.I(\mod.cpu.bufreg2.i_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__I0 (.I(\mod.cpu.bufreg2.i_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(\mod.cpu.bufreg2.i_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A1 (.I(\mod.cpu.bufreg2.i_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__I0 (.I(\mod.cpu.bufreg2.i_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(\mod.cpu.bufreg2.i_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A1 (.I(\mod.cpu.bufreg2.i_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__I0 (.I(\mod.cpu.bufreg2.i_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__I1 (.I(\mod.cpu.bufreg2.i_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A1 (.I(\mod.cpu.bufreg2.i_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__I0 (.I(\mod.cpu.bufreg2.i_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__I1 (.I(\mod.cpu.bufreg2.i_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(\mod.cpu.bufreg2.i_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__A1 (.I(\mod.cpu.bufreg2.i_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(\mod.cpu.bufreg2.i_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A1 (.I(\mod.cpu.bufreg2.i_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A1 (.I(\mod.cpu.bufreg2.i_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(\mod.cpu.bufreg2.i_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1154__I (.I(\mod.cpu.bufreg2.i_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(\mod.cpu.bufreg2.i_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1503__I (.I(\mod.cpu.bufreg2.i_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(\mod.cpu.bufreg2.i_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__I (.I(\mod.cpu.bufreg2.i_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1118__I (.I(\mod.cpu.bufreg2.i_op_b_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__A1 (.I(\mod.cpu.bufreg2.i_op_b_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1017__I (.I(\mod.cpu.bufreg2.i_op_b_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__A1 (.I(\mod.cpu.bufreg2.i_op_b_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1103__A1 (.I(\mod.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1071__I (.I(\mod.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A3 (.I(\mod.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__A1 (.I(\mod.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__B2 (.I(\mod.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__A1 (.I(\mod.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A1 (.I(\mod.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1120__B1 (.I(\mod.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1112__I (.I(\mod.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1101__I (.I(\mod.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1021__A1 (.I(\mod.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1018__A1 (.I(\mod.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__B1 (.I(\mod.cpu.i_rf_ready ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1044__I0 (.I(\mod.cpu.i_rf_ready ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__I0 (.I(\mod.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__I1 (.I(\mod.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1158__A4 (.I(\mod.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1019__A2 (.I(\mod.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(\mod.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__I1 (.I(\mod.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__I1 (.I(\mod.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1158__A1 (.I(\mod.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(\mod.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A1 (.I(\mod.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__I1 (.I(\mod.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1161__A1 (.I(\mod.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A2 (.I(\mod.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__I1 (.I(\mod.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1037__I1 (.I(\mod.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__B (.I(\mod.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A1 (.I(\mod.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(\mod.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__I1 (.I(\mod.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A1 (.I(\mod.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__I1 (.I(\mod.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A1 (.I(\mod.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A1 (.I(\mod.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__I0 (.I(\mod.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__C (.I(\mod.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1135__I (.I(\mod.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1125__A1 (.I(\mod.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__A1 (.I(\mod.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__A2 (.I(\mod.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A1 (.I(\mod.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__A1 (.I(\mod.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__A1 (.I(\mod.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__D (.I(\mod.u_scanchain_local.module_data_in[95] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1060__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__CLKN (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1043 ();
 assign io_oeb[0] = net8;
 assign io_oeb[10] = net18;
 assign io_oeb[11] = net19;
 assign io_oeb[12] = net20;
 assign io_oeb[13] = net21;
 assign io_oeb[14] = net22;
 assign io_oeb[15] = net23;
 assign io_oeb[16] = net24;
 assign io_oeb[17] = net25;
 assign io_oeb[18] = net26;
 assign io_oeb[19] = net27;
 assign io_oeb[1] = net9;
 assign io_oeb[20] = net28;
 assign io_oeb[21] = net29;
 assign io_oeb[22] = net30;
 assign io_oeb[23] = net31;
 assign io_oeb[24] = net32;
 assign io_oeb[25] = net33;
 assign io_oeb[26] = net34;
 assign io_oeb[27] = net35;
 assign io_oeb[28] = net36;
 assign io_oeb[29] = net37;
 assign io_oeb[2] = net10;
 assign io_oeb[30] = net38;
 assign io_oeb[31] = net39;
 assign io_oeb[32] = net40;
 assign io_oeb[33] = net41;
 assign io_oeb[34] = net42;
 assign io_oeb[35] = net43;
 assign io_oeb[36] = net44;
 assign io_oeb[37] = net45;
 assign io_oeb[3] = net11;
 assign io_oeb[4] = net12;
 assign io_oeb[5] = net13;
 assign io_oeb[6] = net14;
 assign io_oeb[7] = net15;
 assign io_oeb[8] = net16;
 assign io_oeb[9] = net17;
 assign io_out[0] = net46;
 assign io_out[10] = net56;
 assign io_out[11] = net57;
 assign io_out[12] = net58;
 assign io_out[13] = net59;
 assign io_out[14] = net60;
 assign io_out[15] = net61;
 assign io_out[19] = net62;
 assign io_out[1] = net47;
 assign io_out[20] = net63;
 assign io_out[21] = net64;
 assign io_out[22] = net65;
 assign io_out[23] = net66;
 assign io_out[24] = net67;
 assign io_out[25] = net68;
 assign io_out[26] = net69;
 assign io_out[27] = net70;
 assign io_out[28] = net71;
 assign io_out[29] = net72;
 assign io_out[2] = net48;
 assign io_out[30] = net73;
 assign io_out[31] = net74;
 assign io_out[32] = net75;
 assign io_out[33] = net76;
 assign io_out[34] = net77;
 assign io_out[35] = net78;
 assign io_out[36] = net79;
 assign io_out[37] = net80;
 assign io_out[3] = net49;
 assign io_out[4] = net50;
 assign io_out[5] = net51;
 assign io_out[6] = net52;
 assign io_out[7] = net53;
 assign io_out[8] = net54;
 assign io_out[9] = net55;
 assign la_data_out[0] = net81;
 assign la_data_out[10] = net91;
 assign la_data_out[11] = net92;
 assign la_data_out[12] = net93;
 assign la_data_out[13] = net94;
 assign la_data_out[14] = net95;
 assign la_data_out[15] = net96;
 assign la_data_out[16] = net97;
 assign la_data_out[17] = net98;
 assign la_data_out[18] = net99;
 assign la_data_out[19] = net100;
 assign la_data_out[1] = net82;
 assign la_data_out[20] = net101;
 assign la_data_out[21] = net102;
 assign la_data_out[22] = net103;
 assign la_data_out[23] = net104;
 assign la_data_out[24] = net105;
 assign la_data_out[25] = net106;
 assign la_data_out[26] = net107;
 assign la_data_out[27] = net108;
 assign la_data_out[28] = net109;
 assign la_data_out[29] = net110;
 assign la_data_out[2] = net83;
 assign la_data_out[30] = net111;
 assign la_data_out[31] = net112;
 assign la_data_out[32] = net113;
 assign la_data_out[33] = net114;
 assign la_data_out[34] = net115;
 assign la_data_out[35] = net116;
 assign la_data_out[36] = net117;
 assign la_data_out[37] = net118;
 assign la_data_out[38] = net119;
 assign la_data_out[39] = net120;
 assign la_data_out[3] = net84;
 assign la_data_out[40] = net121;
 assign la_data_out[41] = net122;
 assign la_data_out[42] = net123;
 assign la_data_out[43] = net124;
 assign la_data_out[44] = net125;
 assign la_data_out[45] = net126;
 assign la_data_out[46] = net127;
 assign la_data_out[47] = net128;
 assign la_data_out[48] = net129;
 assign la_data_out[49] = net130;
 assign la_data_out[4] = net85;
 assign la_data_out[50] = net131;
 assign la_data_out[51] = net132;
 assign la_data_out[52] = net133;
 assign la_data_out[53] = net134;
 assign la_data_out[54] = net135;
 assign la_data_out[55] = net136;
 assign la_data_out[56] = net137;
 assign la_data_out[57] = net138;
 assign la_data_out[58] = net139;
 assign la_data_out[59] = net140;
 assign la_data_out[5] = net86;
 assign la_data_out[60] = net141;
 assign la_data_out[61] = net142;
 assign la_data_out[62] = net143;
 assign la_data_out[63] = net144;
 assign la_data_out[6] = net87;
 assign la_data_out[7] = net88;
 assign la_data_out[8] = net89;
 assign la_data_out[9] = net90;
 assign user_irq[0] = net145;
 assign user_irq[1] = net146;
 assign user_irq[2] = net147;
 assign wbs_ack_o = net148;
 assign wbs_dat_o[0] = net149;
 assign wbs_dat_o[10] = net159;
 assign wbs_dat_o[11] = net160;
 assign wbs_dat_o[12] = net161;
 assign wbs_dat_o[13] = net162;
 assign wbs_dat_o[14] = net163;
 assign wbs_dat_o[15] = net164;
 assign wbs_dat_o[16] = net165;
 assign wbs_dat_o[17] = net166;
 assign wbs_dat_o[18] = net167;
 assign wbs_dat_o[19] = net168;
 assign wbs_dat_o[1] = net150;
 assign wbs_dat_o[20] = net169;
 assign wbs_dat_o[21] = net170;
 assign wbs_dat_o[22] = net171;
 assign wbs_dat_o[23] = net172;
 assign wbs_dat_o[24] = net173;
 assign wbs_dat_o[25] = net174;
 assign wbs_dat_o[26] = net175;
 assign wbs_dat_o[27] = net176;
 assign wbs_dat_o[28] = net177;
 assign wbs_dat_o[29] = net178;
 assign wbs_dat_o[2] = net151;
 assign wbs_dat_o[30] = net179;
 assign wbs_dat_o[31] = net180;
 assign wbs_dat_o[3] = net152;
 assign wbs_dat_o[4] = net153;
 assign wbs_dat_o[5] = net154;
 assign wbs_dat_o[6] = net155;
 assign wbs_dat_o[7] = net156;
 assign wbs_dat_o[8] = net157;
 assign wbs_dat_o[9] = net158;
endmodule

