* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_ip_sram__sram256x8m8wm1 abstract view
.subckt gf180mcu_fd_ip_sram__sram256x8m8wm1 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7]
+ CEN CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] GWEN Q[0] Q[1] Q[2] Q[3] Q[4] Q[5]
+ Q[6] Q[7] WEN[0] WEN[1] WEN[2] WEN[3] WEN[4] WEN[5] WEN[6] WEN[7] VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA_mod.u_scanchain_local.scan_flop\[57\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2479__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2106_ _0464_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3086_ la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _0424_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _2939_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_85_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1445__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1996__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[3\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2173__A2 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1684__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1389__I _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1987__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ _0133_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ _0068_ io_in[12] mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1606_ _1043_ _1048_ mod.u_arbiter.o_wb_cpu_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2013__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2586_ _0012_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1537_ mod.u_cpu.cpu.decode.op21 _0829_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1372__B1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1468_ _0922_ mod.u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1399_ _0857_ _0868_ _0881_ mod.u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_cpu.rf_ram.RAM0_GWEN _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[15\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1363__B1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1666__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2672__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_mod.u_scanchain_local.scan_flop\[22\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1969__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2440_ _0241_ _0384_ _0534_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2371_ _0521_ _0680_ _0681_ _1156_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[38\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2452__B _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _0116_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2385__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ _0051_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2569_ _0928_ _0267_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2695__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1515__C _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1648__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2119__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2346__C _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1757__I _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1820__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1423__I1 mod.u_cpu.rf_ram.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2376__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2533__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1351__A3 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1639__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1940_ _0323_ _0251_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1871_ _0285_ _0278_ _0287_ _1030_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2423_ _0834_ _0390_ _0649_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2354_ _0371_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2285_ _0400_ _0337_ _0532_ _0603_ _0368_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2447__B _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2515__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2294__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2710__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[49\] mod.u_scanchain_local.module_data_in\[48\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[11\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_54_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2972_ io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _0310_ _0321_ _0311_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1854_ _0272_ mod.u_cpu.cpu.genblk3.csr.mcause31 _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1785_ mod.u_cpu.rf_ram_if.rcnt\[0\] _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2406_ _0256_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2337_ mod.u_cpu.cpu.immdec.imm30_25\[3\] _0390_ _0635_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2268_ _0584_ _0587_ _0588_ _0568_ _0408_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2276__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2733__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2276__B2 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2199_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2028__B2 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2503__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2267__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2019__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _0859_ _1016_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2606__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1881__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2756__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _0474_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _0432_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2258__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2886_ _2886_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1906_ _1046_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2430__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2460__B _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1837_ _0938_ _0846_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1768_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2194__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _1053_ _1117_ _1118_ mod.u_arbiter.o_wb_cpu_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2497__A1 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2249__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2127__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2629__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2421__A1 mod.u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2779__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1932__B1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ _0149_ io_in[12] mod.u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2412__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2671_ _0083_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1766__A3 mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ _1038_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1553_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1484_ _0926_ _0931_ _0932_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2479__A1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2479__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2105_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] _1143_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3085_ la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2036_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\]
+ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2938_ _2938_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2403__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2190__B _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _2869_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2621__D _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[3\]_D mod.u_arbiter.i_wb_cpu_rdt\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1445__A2 _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[31\] mod.u_arbiter.i_wb_cpu_rdt\[28\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2330__B1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2723_ _0132_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2654_ _0067_ io_in[12] mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1605_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1046_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2585_ _0011_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1536_ _0842_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1372__A1 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1372__B2 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1467_ mod.u_cpu.rf_ram_if.wdata0_r\[3\] mod.u_cpu.rf_ram_if.wdata1_r\[3\] _0865_
+ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1398_ _0868_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2172__I0 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3068_ la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2019_ _0390_ _0311_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__B1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1363__B2 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1910__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2095__B _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_scanchain_local.scan_flop\[41\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2091__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[56\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ _0940_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_mod.u_scanchain_local.clk mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2082__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2452__C _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _0115_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2637_ _0050_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2542__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2568_ _0928_ _0267_ _0819_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2499_ mod.u_arbiter.i_wb_cpu_rdt\[10\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _0750_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1519_ _0933_ _0941_ _0945_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[3\] mod.u_arbiter.i_wb_cpu_rdt\[0\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ clknet_3_0__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2135__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1820__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1959__I0 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1584__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2533__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1811__A2 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1870_ _0286_ _0844_ _0278_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2422_ _0715_ _0687_ _0720_ _0727_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2353_ _0339_ _0357_ _0665_ _0252_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2127__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2284_ _0379_ _0527_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1999_ _0245_ _0252_ _0355_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2662__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__B _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[12\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2515__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2515__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2294__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2046__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2109__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[28\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2285__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1879__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2971_ io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ _0319_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2685__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1853_ _0846_ _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1548__A1 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1784_ mod.u_cpu.rf_ram_if.rcnt\[0\] _0823_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _0325_ _0711_ _0675_ _0339_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1720__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2336_ _0639_ _0637_ _0649_ _0650_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2267_ _0251_ _0335_ _0579_ _0252_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ _0958_ _0523_ _0218_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2028__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2193__B _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2413__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2200__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[61\] mod.u_scanchain_local.module_data_in\[60\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[23\] clknet_3_2__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2019__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1950__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] mod.u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _1164_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2052_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\]
+ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2954_ _2954_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1769__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2885_ _2885_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1905_ mod.u_arbiter.i_wb_cpu_ack mod.u_arbiter.o_wb_cpu_adr\[1\] _0305_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2430__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1836_ _0256_ _0260_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1767_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1698_ mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] _1073_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1941__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2700__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2497__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2319_ _0258_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2619__D _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2249__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2421__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2143__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2185__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1932__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1730__B _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2670_ _0082_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2280__C _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1621_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _1056_
+ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2723__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1923__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[18\]_D mod.u_arbiter.i_wb_cpu_rdt\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1552_ mod.u_cpu.cpu.state.o_cnt_r\[2\] mod.u_cpu.cpu.ctrl.i_iscomp _0929_ _1002_
+ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1483_ _0828_ _0933_ mod.u_cpu.cpu.decode.co_ebreak _0829_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2479__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2104_ _1143_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3084_ la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_78_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2035_ _0423_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2100__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2937_ _2937_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2471__B mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2403__A2 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2868_ _2868_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2167__A1 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2799_ _0208_ io_in[12] mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1819_ _0242_ _0243_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1914__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[24\] mod.u_arbiter.i_wb_cpu_rdt\[21\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2746__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1905__A1 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__B2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1887__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2722_ _0131_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2397__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2397__B2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2653_ _0066_ io_in[12] mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1604_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1046_ _1041_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2584_ _0010_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1535_ _0968_ _0969_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1372__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1466_ _0921_ mod.u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2321__A1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1397_ _0865_ _0878_ _0859_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2619__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2172__I1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3067_ la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2018_ _0255_ _0380_ _0385_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2769__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2388__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1363__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[61\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2163__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2312__B2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2312__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1666__A3 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__I1 mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2076__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2379__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2551__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0114_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _0049_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2542__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2567_ _0928_ _0267_ _1036_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2542__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2498_ _0781_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1518_ _0967_ mod.u_cpu.rf_ram_if.rdata1\[0\] _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1449_ mod.u_cpu.rf_ram_if.rdata1\[1\] _0895_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3119_ wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_93_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2151__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1584__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A1 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1895__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2553__C _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1811__A3 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2421_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _0376_ _0723_ _0726_ _0687_ _0727_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2352_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_arbiter.i_wb_cpu_rdt\[12\] _1046_ _0665_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2283_ _0593_ _0525_ _0601_ _0602_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1998_ _0371_ _0391_ _0393_ _0368_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2619_ _0020_ io_in[12] mod.u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_mod.u_scanchain_local.scan_flop\[40\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[55\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1895__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[12\] _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2293__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1852_ _0944_ mod.u_cpu.cpu.decode.co_ebreak _0832_ _0988_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1783_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r mod.u_cpu.cpu.state.stage_two_req
+ _0218_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1548__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2404_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2335_ mod.u_cpu.cpu.immdec.imm30_25\[2\] _0634_ _0376_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1720__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2266_ _0247_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2197_ _0939_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1484__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1869__I mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[54\] mod.u_scanchain_local.module_data_in\[53\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[16\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_72_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1728__B _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[6\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2120_ _0473_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2051_ _0431_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2652__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2953_ _2953_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1904_ _0304_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _2884_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ mod.u_cpu.cpu.ctrl.i_iscomp _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1766_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] mod.u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2194__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1941__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2318_ _0958_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2249_ _0330_ _0365_ _0349_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1599__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[18\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2185__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1932__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2675__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1999__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1471__I1 mod.u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1620_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _1056_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\]
+ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1551_ _1001_ mod.u_cpu.cpu.ctrl.i_iscomp _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1923__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1482_ mod.u_arbiter.i_wb_cpu_dbus_we _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2103_ _1159_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3083_ la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2034_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2936_ _2936_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2867_ _2867_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1818_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[0\] _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2167__A2 mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2798_ _0207_ io_in[12] mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ _0827_ mod.u_cpu.cpu.decode.opcode\[1\] _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2698__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1914__A2 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[17\] mod.u_arbiter.i_wb_cpu_rdt\[14\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2721_ _0130_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2397__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ _0065_ io_in[12] mod.u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1603_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2583_ _0009_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1534_ _0974_ _0979_ _0983_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1465_ mod.u_cpu.rf_ram_if.wdata0_r\[2\] mod.u_cpu.rf_ram_if.wdata1_r\[2\] _0865_
+ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1396_ mod.u_cpu.cpu.decode.op26 mod.u_cpu.cpu.decode.co_ebreak _0865_ _0879_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2321__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3066_ la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2017_ _0244_ _0249_ _0379_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2919_ _2919_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__A2 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2149__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2312__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2713__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2567__B _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1814__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2704_ _0113_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ _0048_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2527__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2542__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2566_ _1035_ _0267_ _0818_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2497_ mod.u_arbiter.i_wb_cpu_rdt\[9\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] _0750_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1517_ mod.u_cpu.rf_ram.regzero _0967_ _0888_ _0890_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1448_ mod.u_cpu.rf_ram_if.rtrig1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2736__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3118_ wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1379_ mod.u_cpu.rf_ram_if.wen1_r _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3049_ la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2230__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2297__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2609__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2509__C1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1980__B1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0364_ _0724_ _0725_ _0253_ _0256_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2351_ _0366_ _0625_ _0662_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2759__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2282_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _0376_ _0525_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2288__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1421__S mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2460__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1997_ _0352_ _0365_ _0392_ _0357_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2212__B2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[51\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ _0019_ io_in[12] mod.u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2549_ _0807_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2515__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2279__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2203__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1920_ _1045_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2293__I1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2442__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1851_ _0952_ _1030_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1782_ _0217_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1548__A3 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2581__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ _1046_ mod.u_arbiter.i_wb_cpu_rdt\[23\] _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2334_ _0308_ _0640_ _0648_ _0409_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2265_ _0253_ _0325_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2196_ _0826_ _0926_ _0931_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2157__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[47\] mod.u_scanchain_local.module_data_in\[46\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[9\] clknet_3_4__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2424__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1744__B _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2050_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\]
+ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2952_ _2952_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2415__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1903_ mod.u_arbiter.i_wb_cpu_rdt\[31\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _0288_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2883_ _2883_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1834_ _0258_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_mod.u_scanchain_local.scan_flop\[54\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1765_ _0957_ _1142_ _0949_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1696_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] _1111_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[69\]_CLK clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2317_ _0926_ _0933_ _1144_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2248_ _0245_ _0325_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_39_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2179_ _0500_ _0505_ _0507_ _0973_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2406__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1829__B _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1393__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[6\]_D mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__A3 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1739__B _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_67_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1384__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1481_ _0926_ mod.u_cpu.cpu.decode.opcode\[1\] _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1687__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2102_ _0826_ _0946_ _1161_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3082_ la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2033_ _0422_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_36_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _2935_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2866_ _2866_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1817_ _1045_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2167__A3 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2797_ _0206_ io_in[12] mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1748_ _1151_ _1154_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1679_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _1100_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2642__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1669__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2792__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1841__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ _0129_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2651_ _0064_ io_in[12] mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1602_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2582_ _0008_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1533_ _0826_ _0955_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1464_ _0920_ mod.u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1395_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3065_ la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2016_ _0259_ _0400_ _0401_ _0410_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_36_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1832__A2 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _2918_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2665__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2849_ _2849_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_12_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1520__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2076__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2165__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1823__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1511__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2688__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1578__A1 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2703_ _0112_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2634_ _0047_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2565_ mod.u_cpu.cpu.state.o_cnt_r\[3\] mod.u_cpu.cpu.state.o_cnt\[2\] _0818_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2527__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2527__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1516_ _0912_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2496_ _0780_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1750__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1447_ _0911_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1378_ mod.u_cpu.rf_ram_if.genblk1.wtrig0_r _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3117_ wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_71_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3048_ la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1569__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2230__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1741__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2509__C2 mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2509__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1980__B2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1732__A1 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ _0334_ _0357_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2281_ _0390_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2288__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1501__I mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _0334_ _0365_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1971__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2703__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ _0018_ io_in[12] mod.u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2548_ mod.u_cpu.cpu.state.o_cnt\[2\] _0928_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0210_
+ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1574__I1 mod.u_cpu.rf_ram.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1392__B _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2479_ mod.u_arbiter.i_wb_cpu_rdt\[3\] _0744_ _0750_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2279__A2 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1411__I mod.u_cpu.rf_ram.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[1\] mod.timer_irq io_in[11] mod.u_arbiter.o_wb_cpu_we
+ clknet_3_3__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_54_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1567__B _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2203__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1962__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2442__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _0996_ _0261_ _0271_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1781_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _0215_ _0216_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1548__A4 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1953__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2402_ _0544_ _0626_ _0707_ _0708_ _0693_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_44_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1705__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ _0364_ _0641_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_3__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2264_ _0335_ _0569_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2195_ mod.u_cpu.cpu.immdec.imm19_12_20\[0\] _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ _0258_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2749__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2188__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1935__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2360__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1760__B _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[41\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2951_ _2951_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ _0303_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2882_ _2882_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1833_ mod.u_arbiter.i_wb_cpu_ack _1038_ _0257_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1764_ _1053_ _1167_ mod.u_arbiter.o_wb_cpu_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1926__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1695_ _1053_ _1114_ _1115_ mod.u_arbiter.o_wb_cpu_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2316_ _0621_ _0622_ _0218_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ _0249_ _0332_ _0355_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_39_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2178_ _0506_ _0930_ _0500_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2342__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[64\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2030__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1908__A1 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ _0825_ mod.u_cpu.cpu.decode.opcode\[1\] _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2333__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ _1139_ _0460_ _0461_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3081_ la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2032_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2934_ _2934_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2865_ _2865_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1816_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2796_ _0205_ io_in[12] mod.u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1747_ mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1152_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2572__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1678_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _1100_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2088__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1366__A2 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2315__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[53\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2094__A3 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[68\]_CLK clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2650_ _0063_ io_in[12] mod.u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ mod.u_cpu.cpu.genblk1.align.ctrl_misal _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2581_ _0007_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1532_ _0980_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1463_ mod.u_cpu.rf_ram_if.wdata0_r\[1\] mod.u_cpu.rf_ram_if.wdata1_r\[1\] _0865_
+ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2157__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2306__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1932__C _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1394_ _0861_ _0868_ _0877_ mod.u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3064_ la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2015_ _0376_ _0403_ _0406_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2917_ _2917_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1596__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2848_ _2848_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2779_ _0188_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2545__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1520__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2245__I mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2233__B1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[22\] mod.u_arbiter.i_wb_cpu_rdt\[19\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0111_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1994__I _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2633_ _0046_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2527__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2564_ _1035_ _1001_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1515_ mod.u_arbiter.i_wb_cpu_dbus_we mod.u_cpu.cpu.bufreg.i_sh_signed _0831_ _0827_
+ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1943__B _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2495_ mod.u_arbiter.i_wb_cpu_rdt\[8\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] _0750_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1446_ mod.u_cpu.rf_ram_if.rdata0\[7\] _0910_ mod.u_cpu.rf_ram_if.rtrig0 _0911_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1377_ _0863_ _0864_ mod.u_arbiter.i_wb_cpu_dbus_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1502__A2 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3116_ wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3047_ la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2463__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2632__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2782__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[9\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A1 mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2509__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1732__A2 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _0364_ _0596_ _0597_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2655__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__B1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _0249_ _0352_ _0357_ _0252_ _0365_ _0314_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1420__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2616_ _0017_ io_in[12] mod.u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1971__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2547_ _0806_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2478_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _1168_ _0757_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1429_ _0900_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1962__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1602__I _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1780_ mod.u_arbiter.i_wb_cpu_ack _1038_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1402__B2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1953__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2401_ _0241_ _0336_ _0313_ _0244_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2332_ _0247_ _0643_ _0646_ _0517_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2263_ _0335_ _0340_ _0341_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2194_ _0511_ _0259_ _0518_ _0520_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__B1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ _0874_ _0346_ _0374_ _0375_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1632__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2188__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1935__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1699__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2360__A2 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _2950_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_90_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2881_ _2881_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1901_ mod.u_arbiter.i_wb_cpu_rdt\[30\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0288_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1832_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _0215_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1763_ mod.u_cpu.cpu.state.init_done _0990_ _1144_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] _1073_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1926__A2 mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2315_ _0332_ _0371_ _0629_ _0630_ _0255_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1443__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2246_ _0339_ _0371_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2177_ mod.u_cpu.cpu.alu.cmp_r _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1862__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1862__B2 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1917__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__B _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2716__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[52\] mod.u_scanchain_local.module_data_in\[51\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[14\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_60_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1369__B1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2030__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1908__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__B _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _0864_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3080_ la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _0421_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_48_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1844__A1 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2933_ _2933_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_51_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2864_ _2864_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_141_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1815_ _1045_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2795_ _0204_ io_in[12] mod.u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1438__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1746_ _0937_ _0962_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2572__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1677_ _1042_ _1100_ _1101_ _1102_ mod.u_arbiter.o_wb_cpu_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2739__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1901__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ mod.u_cpu.cpu.immdec.imm19_12_20\[2\] _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__A1 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1438__I1 mod.u_cpu.rf_ram.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[31\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1366__A3 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1600_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2539__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2003__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2580_ _0006_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1762__B1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1531_ _0830_ _0839_ mod.u_cpu.cpu.alu.cmp_r _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1462_ _0919_ mod.u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2306__A2 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1393_ _0865_ _0875_ _0876_ _0868_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3063_ la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1817__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ _0258_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_1_0_mod.u_scanchain_local.clk clknet_3_2__leaf_mod.u_scanchain_local.clk
+ clknet_opt_1_0_mod.u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2916_ _2916_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2242__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ _2847_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_mod.u_scanchain_local.scan_flop\[54\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2778_ _0187_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1729_ _1139_ _0864_ _0837_ mod.u_arbiter.i_wb_cpu_dbus_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2545__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__A3 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1808__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2481__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2233__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xmod.u_scanchain_local.scan_flop\[15\] mod.u_arbiter.i_wb_cpu_rdt\[12\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] clknet_3_0__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2210__B _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2472__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2224__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2224__B2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2701_ _0110_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1496__B mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2584__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _0045_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2527__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2563_ _0817_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1514_ mod.u_cpu.cpu.alu.add_cy_r mod.u_cpu.cpu.alu.i_rs1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2494_ _0779_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1445_ _0887_ _0023_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1376_ mod.u_cpu.cpu.bufreg.lsb\[0\] _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1502__A3 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3115_ wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1451__S _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3046_ la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__B1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[52\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[67\]_CLK clknet_3_2__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2256__I mod.u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2192__S _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2206__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2509__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1335__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1496__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__B2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _0218_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1420__A2 _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ _0025_ io_in[12] mod.u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1559__I0 mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1446__S mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ _1036_ mod.u_cpu.cpu.state.o_cnt_r\[2\] _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ _1168_ _1170_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1428_ mod.u_cpu.rf_ram.rdata\[3\] mod.u_cpu.rf_ram.data\[3\] _0026_ _0900_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1359_ _0833_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3029_ la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2436__A1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1478__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2427__A1 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1650__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1402__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2400_ _0317_ _0404_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2622__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2331_ _0625_ _0644_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2262_ _0340_ _0512_ _0581_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_78_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2772__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ _0408_ _0519_ _0376_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2418__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2418__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _0259_ _0346_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2529_ mod.u_arbiter.i_wb_cpu_rdt\[25\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] _0777_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[6\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2188__A3 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[9\]_D mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2795__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1623__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1900_ _0302_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0218_ _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1762_ _0830_ _0863_ _0864_ _0831_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1693_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] _1111_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_100_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2336__B1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2314_ _0244_ _0514_ _0371_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ mod.u_cpu.cpu.csr_imm _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2176_ _1033_ _0503_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1862__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1614__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__B _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.output_buffers\[2\]_I mod.u_scanchain_local.data_out_i
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[45\] mod.u_scanchain_local.module_data_in\[44\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[7\] clknet_3_4__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1605__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1369__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2030__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2169__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1541__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2097__A2 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2932_ _2932_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2863_ _2863_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2794_ _0203_ io_in[12] mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1814_ _1035_ _0239_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1745_ _0936_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2021__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2572__A3 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1676_ mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] _1041_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1780__A1 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2088__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2228_ _0542_ _0525_ _0551_ _0552_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2159_ mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] mod.u_arbiter.i_wb_cpu_dbus_adr\[28\]
+ _1163_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1835__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1771__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_mod.u_scanchain_local.clk_I mod.u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2251__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2539__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2539__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2003__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1762__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1530_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _0929_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1762__B2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1461_ mod.u_cpu.rf_ram_if.wdata0_r\[0\] mod.u_cpu.rf_ram_if.wdata1_r\[0\] _0865_
+ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1392_ _0835_ _0846_ _0865_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3062_ la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1817__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ _2915_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1449__S _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2242__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2846_ _2846_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2706__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2777_ _0186_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1728_ _1139_ _1140_ _0837_ mod.u_arbiter.i_wb_cpu_dbus_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1659_ _1042_ _1087_ _1088_ _1089_ mod.u_arbiter.o_wb_cpu_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_63_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1505__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1912__S _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2233__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[11\]_D mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2224__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0109_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2729__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1983__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2631_ _0044_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ _1036_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1513_ _0930_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2401__B _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2493_ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] _0757_ _0777_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ mod.u_arbiter.i_wb_cpu_rdt\[7\] _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1444_ _0909_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1375_ mod.u_cpu.cpu.bufreg.lsb\[1\] _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1502__A4 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3114_ wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3045_ la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[21\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2215__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1974__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2829_ _2829_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__1974__B2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2311__B _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1965__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1717__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2390__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[44\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2594__D mod.u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__A2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _0346_ _0377_ _0378_ _0389_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0036_ io_in[12] mod.u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1708__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1559__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0938_ _1143_ _0805_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2381__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2476_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _1169_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1427_ _0899_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1358_ _0842_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3028_ io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2293__S _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2306__B _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1947__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[67\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1478__A3 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2574__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2427__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2060__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1938__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2363__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _0334_ _0349_ _0365_ _0544_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2261_ _0323_ _0379_ _0335_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2192_ mod.u_arbiter.i_wb_cpu_rdt\[31\] mod.u_arbiter.i_wb_cpu_rdt\[15\] _1046_ _0519_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2418__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[51\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1976_ _0308_ _0349_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_mod.u_scanchain_local.scan_flop\[66\]_CLK clknet_3_2__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1929__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1457__S _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2354__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2528_ _0796_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[19\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2188__A4 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__A2 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2345__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ _0245_ _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1761_ _0933_ _1038_ mod.u_arbiter.o_wb_cpu_we vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1692_ _1042_ _1111_ _1112_ _1113_ mod.u_arbiter.o_wb_cpu_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2313_ _0625_ _0628_ _0342_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2244_ _0561_ _0525_ _0565_ _0566_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2175_ mod.u_cpu.cpu.alu.i_rs1 _0502_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1959_ mod.u_arbiter.i_wb_cpu_rdt\[9\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _1044_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1915__S _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2327__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2327__B2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2612__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[38\] mod.u_scanchain_local.module_data_in\[37\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[0\] clknet_3_3__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2566__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2015__B1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1369__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2762__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1825__S _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2318__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_cpu.rf_ram.RAM0 mod.u_cpu.rf_ram.RAM0/A[0] mod.u_cpu.rf_ram.RAM0/A[1] mod.u_cpu.rf_ram.RAM0/A[2]
+ mod.u_cpu.rf_ram.RAM0/A[3] mod.u_cpu.rf_ram.RAM0/A[4] mod.u_cpu.rf_ram.RAM0/A[5]
+ mod.u_cpu.rf_ram.RAM0/A[6] mod.u_cpu.rf_ram.RAM0/A[7] mod.u_cpu.rf_ram.RAM0/CEN
+ mod.u_cpu.rf_ram.RAM0/CLK mod.u_cpu.rf_ram.RAM0/D[0] mod.u_cpu.rf_ram.RAM0/D[1]
+ mod.u_cpu.rf_ram.RAM0/D[2] mod.u_cpu.rf_ram.RAM0/D[3] mod.u_cpu.rf_ram.RAM0/D[4]
+ mod.u_cpu.rf_ram.RAM0/D[5] mod.u_cpu.rf_ram.RAM0/D[6] mod.u_cpu.rf_ram.RAM0/D[7]
+ mod.u_cpu.rf_ram.RAM0/GWEN mod.u_cpu.rf_ram.RAM0/Q[0] mod.u_cpu.rf_ram.RAM0/Q[1]
+ mod.u_cpu.rf_ram.RAM0/Q[2] mod.u_cpu.rf_ram.RAM0/Q[3] mod.u_cpu.rf_ram.RAM0/Q[4]
+ mod.u_cpu.rf_ram.RAM0/Q[5] mod.u_cpu.rf_ram.RAM0/Q[6] mod.u_cpu.rf_ram.RAM0/Q[7]
+ mod.u_cpu.rf_ram.RAM0/WEN[0] mod.u_cpu.rf_ram.RAM0/WEN[1] mod.u_cpu.rf_ram.RAM0/WEN[2]
+ mod.u_cpu.rf_ram.RAM0/WEN[3] mod.u_cpu.rf_ram.RAM0/WEN[4] mod.u_cpu.rf_ram.RAM0/WEN[5]
+ mod.u_cpu.rf_ram.RAM0/WEN[6] mod.u_cpu.rf_ram.RAM0/WEN[7] vdd vss gf180mcu_fd_ip_sram__sram256x8m8wm1
XFILLER_36_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2931_ _2931_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2254__B1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2391__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2862_ _2862_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2793_ _0202_ io_in[12] mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1813_ _0944_ mod.u_cpu.cpu.genblk3.csr.o_new_irq _0235_ _0238_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2557__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1744_ _1149_ _1150_ _1151_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1675_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _1096_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1780__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ mod.u_cpu.cpu.immdec.imm19_12_20\[2\] _0259_ _0525_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _0492_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2493__C2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2493__B1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2635__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2089_ _0451_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_scanchain_local.input_buf_clk_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2785__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__B _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2484__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1995__C1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2539__A1 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2539__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2003__A3 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1762__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1460_ _0918_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1354__I mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1391_ _0874_ _0859_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3130_ mod.u_scanchain_local.data_out io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1514__A2 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3061_ la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2012_ _0245_ _0254_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2914_ _2914_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1825__I0 mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2845_ _2845_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2776_ _0185_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1727_ mod.u_cpu.cpu.bne_or_bge _0864_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1465__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1658_ mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] _1073_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1505__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1589_ _0990_ _1033_ _1034_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2800__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1349__I mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1983__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ _0043_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2561_ _1035_ _0816_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2492_ _1177_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1512_ _0937_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1443_ mod.u_cpu.rf_ram.rdata\[6\] mod.u_cpu.rf_ram.data\[6\] _0026_ _0909_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2401__C _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1374_ _0853_ _0862_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3113_ wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3044_ la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2828_ _2828_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2759_ _0168_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2311__C _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1662__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[20\] mod.u_arbiter.i_wb_cpu_rdt\[17\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1965__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1405__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1992_ _0376_ _0387_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_14_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2613_ mod.u_cpu.cpu.o_wdata0 io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1708__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1559__I2 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0938_ mod.u_cpu.cpu.state.init_done _1036_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2381__A2 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2475_ _0764_ _0765_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1426_ mod.u_cpu.rf_ram_if.rdata0\[3\] _0898_ mod.u_cpu.rf_ram_if.rtrig0 _0899_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1357_ _0843_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3027_ io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1947__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2357__C1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2719__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[68\] mod.u_scanchain_local.module_data_in\[67\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[30\] clknet_3_3__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_28_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1828__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1938__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[11\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2363__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ _0528_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2458__I mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2191_ _0513_ _0516_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0256_ _0370_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1929__A2 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__C _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.output_buffers\[3\] clknet_opt_1_1_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.clk_out vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2527_ mod.u_arbiter.i_wb_cpu_rdt\[24\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _0777_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1473__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2458_ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1409_ mod.u_cpu.rf_ram.regzero _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2511__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2389_ mod.u_cpu.cpu.immdec.imm24_20\[2\] _0686_ _0687_ mod.u_cpu.cpu.immdec.imm24_20\[1\]
+ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1865__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[34\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__A3 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2345__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2691__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2227__B _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1760_ _1157_ _1162_ _1165_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1691_ mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] _1041_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2336__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2312_ _0354_ _0626_ _0627_ _0381_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ mod.u_cpu.cpu.csr_imm _0376_ _0525_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2174_ _0501_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2272__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[57\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1958_ _0335_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1889_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _0288_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2327__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1838__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2263__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2015__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2015__B2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[50\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[65\]_CLK clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1829__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _2930_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2254__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2254__B2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ _2861_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2587__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2006__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2792_ _0201_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1812_ _0236_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1743_ _0958_ _1143_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1674_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _1093_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[18\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.out_flop_CLKN clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2226_ _0390_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2157_ mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] mod.u_arbiter.i_wb_cpu_dbus_adr\[27\]
+ _1163_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2493__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2493__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2088_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2548__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2484__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[50\] mod.u_scanchain_local.module_data_in\[49\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[12\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_77_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1995__B1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__C2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2539__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1390_ mod.u_cpu.cpu.immdec.imm11_7\[0\] _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3060_ la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2011_ _0404_ _0368_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2913_ _2913_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2844_ _2844_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2775_ _0184_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1726_ _0863_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1657_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1085_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1545__I mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1588_ _0958_ _0966_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_101_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2602__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2466__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2752__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2209_ _0252_ _0355_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2209__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1680__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2560_ _0944_ mod.u_cpu.cpu.state.o_cnt_r\[3\] _0990_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2625__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2491_ _0749_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1511_ _0946_ _0948_ _0961_ _0927_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1442_ _0908_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2775__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1373_ _0857_ _0858_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3112_ wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3043_ la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2448__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _2827_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2758_ _0167_ io_in[12] mod.u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1709_ _1053_ _1125_ _1126_ mod.u_arbiter.o_wb_cpu_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2689_ _0101_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2439__A1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[9\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2648__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[13\] mod.u_arbiter.i_wb_cpu_rdt\[10\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2798__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ _0252_ _0335_ _0353_ _0249_ _0371_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1405__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2612_ mod.u_cpu.rf_ram_if.wdata0_r\[6\] io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2543_ _0803_ _0804_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1559__I3 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2474_ mod.u_arbiter.i_wb_cpu_rdt\[2\] _0744_ _0750_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1425_ _0887_ _0019_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1356_ mod.u_cpu.cpu.genblk3.csr.o_new_irq _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3026_ io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_93_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2357__B1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1955__I0 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1580__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2060__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ _0321_ _0337_ _0368_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1626__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ _0252_ _0349_ _0354_ _0249_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2423__B _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _0795_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1562__A1 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2457_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1408_ _0851_ _0026_ _0884_ mod.u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2511__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2511__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2388_ _0691_ _0696_ _0390_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1865__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1339_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_72_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3009_ io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2290__A2 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2042__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1608__A2 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2243__B _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1690_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] _1108_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1574__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2311_ _0321_ _0529_ _0527_ _0333_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0376_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2173_ mod.u_cpu.cpu.bne_or_bge mod.u_cpu.cpu.csr_d_sel _0830_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2272__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1957_ _0316_ _0352_ _0353_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_30_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1888_ _0296_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1783__A1 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ mod.u_arbiter.i_wb_cpu_rdt\[15\] _0744_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _0777_ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1535__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2263__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1774__A1 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1829__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2254__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2860_ _2860_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ mod.u_cpu.cpu.genblk3.csr.mie_mtie mod.u_cpu.cpu.genblk3.csr.mstatus_mie mod.timer_irq
+ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2791_ _0200_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2006__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1742_ _1004_ _1005_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ _1053_ _1098_ _1099_ mod.u_arbiter.o_wb_cpu_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2420__C _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2199__I _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ _0368_ _0547_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2156_ _0491_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2493__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[24\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2087_ _0450_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_35_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2548__A3 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2681__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1756__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_mod.u_scanchain_local.scan_flop\[31\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[43\] mod.u_scanchain_local.module_data_in\[42\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[5\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_77_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1995__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1916__I _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_mod.u_scanchain_local.scan_flop\[47\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[14\]_D mod.u_arbiter.i_wb_cpu_rdt\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2010_ _0249_ _0310_ _0364_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_1_0_mod.u_scanchain_local.clk_I clknet_3_2__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2227__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2912_ _2912_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2843_ _2843_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2774_ _0183_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1725_ _1038_ _1137_ _1138_ mod.u_arbiter.o_wb_cpu_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1738__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2431__B _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1656_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1085_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1587_ _0965_ _0972_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2466__A2 mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2208_ _0321_ _0359_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2139_ mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] mod.u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _1163_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A1 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[64\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1729__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2577__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[17\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2209__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ _0776_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1510_ _0864_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1441_ mod.u_cpu.rf_ram_if.rdata0\[6\] _0907_ mod.u_cpu.rf_ram_if.rtrig0 _0908_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3111_ wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1372_ mod.u_cpu.cpu.csr_imm _0824_ _0849_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _0860_
+ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3042_ la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2448__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2826_ _2826_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2757_ _0166_ io_in[12] mod.u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2384__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] _1073_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2688_ _0100_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1639_ _1053_ _1072_ _1074_ mod.u_arbiter.o_wb_cpu_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1505__B _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2439__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2072__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2375__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1990_ _0254_ _0383_ _0386_ _0335_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2611_ mod.u_cpu.rf_ram_if.wdata0_r\[5\] io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2542_ _0501_ _0757_ _0750_ mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] _0804_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2742__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2473_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _1168_ _0757_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1424_ _0897_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1355_ _0826_ _0828_ mod.u_cpu.cpu.decode.op21 _0840_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_96_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3025_ io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2054__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2809_ _2809_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2357__B2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2111__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2615__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1891__I0 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2765__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1399__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2036__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0241_ _0247_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2339__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2525_ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _0757_ _0777_ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ mod.u_arbiter.i_wb_cpu_rdt\[23\] _0778_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1834__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2456_ _1177_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1407_ _0850_ _0868_ _0882_ _0886_ mod.u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2511__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2387_ _0371_ _0382_ _0694_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2638__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1338_ mod.u_cpu.cpu.branch_op _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3008_ io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2788__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1608__A3 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2569__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ _0321_ _0530_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2241_ _0251_ _0408_ _0341_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0946_ _0986_ mod.u_arbiter.i_wb_cpu_dbus_we _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1480__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1956_ mod.u_arbiter.i_wb_cpu_rdt\[2\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _1045_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1887_ mod.u_arbiter.i_wb_cpu_rdt\[23\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _0288_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2508_ _0786_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_1_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1535__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2439_ _0259_ _0734_ _0735_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1774__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2803__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2487__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1810_ _0938_ _1143_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2790_ _0199_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1741_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r _1149_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1672_ mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] _1073_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2224_ _0245_ _0339_ _0548_ _0332_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2429__B _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2155_ mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] mod.u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _1163_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1828__I0 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1939_ _0251_ _0332_ _0334_ _0335_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1756__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2469__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1692__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xmod.u_scanchain_local.scan_flop\[36\] mod.u_scanchain_local.module_data_in\[35\]
+ io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_41_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1995__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2249__B _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _2911_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1435__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1986__A2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2842_ _2842_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2773_ _0182_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1724_ mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] _1038_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1655_ _1042_ _1084_ _1085_ _1086_ mod.u_arbiter.o_wb_cpu_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_mod.u_scanchain_local.scan_flop\[2\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1586_ mod.u_cpu.cpu.alu.add_cy_r mod.u_cpu.cpu.alu.i_rs1 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2207_ _0244_ _0526_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2138_ _0482_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2069_ _0441_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1729__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[14\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2393__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2251__C _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1440_ _0887_ _0022_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1371_ _0835_ _0859_ _0847_ _0824_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3110_ wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3041_ la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2671__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[21\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2825_ _2825_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_143_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2756_ _0165_ io_in[12] mod.u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1707_ _1124_ _1121_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2687_ _0099_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1638_ mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1569_ _0859_ _1017_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1647__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2109__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[8\] mod.u_arbiter.i_wb_cpu_rdt\[5\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ clknet_3_4__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[37\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2694__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1653__A4 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1810__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ mod.u_cpu.rf_ram_if.wdata0_r\[4\] io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2541_ mod.u_arbiter.i_wb_cpu_rdt\[31\] _0744_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2472_ _1168_ _1169_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1423_ mod.u_cpu.rf_ram.rdata\[2\] mod.u_cpu.rf_ram.data\[2\] _0026_ _0897_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1354_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_mod.u_scanchain_local.scan_flop\[63\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1801__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2808_ _2808_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2357__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2739_ _0148_ io_in[12] mod.u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[16\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1891__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2348__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2284__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _0363_ _0364_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_18_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2524_ _0794_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_143_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2455_ _0949_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1406_ mod.u_cpu.cpu.immdec.imm11_7\[4\] _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2386_ _0245_ _0353_ _0527_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2511__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1337_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[66\] mod.u_scanchain_local.module_data_in\[65\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[28\] clknet_3_2__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_56_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2266__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2732__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2018__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2240_ _0318_ _0404_ _0562_ _0530_ _0512_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2171_ _0837_ _0839_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2257__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2009__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ mod.u_arbiter.i_wb_cpu_rdt\[3\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _1045_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1886_ _0295_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2605__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ mod.u_arbiter.i_wb_cpu_rdt\[14\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _0777_ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2438_ mod.u_cpu.cpu.decode.opcode\[1\] _0259_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2369_ _0825_ _0926_ mod.u_cpu.cpu.decode.opcode\[1\] _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2755__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2248__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2117__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__C _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1956__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2420__B2 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2360__B _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2254__C _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2628__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2411__A1 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1740_ _0847_ _0990_ mod.u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1671_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _1096_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2778__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2478__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _0379_ _0368_ _0255_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2154_ _0490_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2085_ _0449_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ _0329_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2402__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1869_ mod.u_cpu.cpu.decode.co_ebreak _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2469__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2469__A1 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[2\]_D mod.u_arbiter.i_wb_cpu_ack vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[29\] mod.u_arbiter.i_wb_cpu_rdt\[26\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_139_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1683__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ _2910_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1435__A2 _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2841_ _2841_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_89_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2772_ _0181_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1723_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1395__I mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] _1073_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1585_ _1030_ _1031_ mod.u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2206_ _0332_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2137_ mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] mod.u_arbiter.i_wb_cpu_dbus_adr\[17\]
+ _1164_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2068_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_4__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1362__A1 mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1665__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2090__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2378__B1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r mod.u_cpu.cpu.genblk3.csr.o_new_irq
+ _0844_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2153__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3040_ la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1408__A2 _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ _2824_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ _0164_ io_in[12] mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1706_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2686_ _0098_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1592__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1637_ _1041_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1568_ _0827_ _0961_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1344__A1 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1499_ mod.u_cpu.cpu.state.stage_two_req _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1647__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2072__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2125__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1583__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1638__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1810__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2540_ _0802_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2471_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] mod.u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1422_ _0896_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2523__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2523__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1353_ _0836_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3023_ io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2054__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ _2807_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_69_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2738_ _0147_ io_in[12] mod.u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2669_ _0081_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1959__S _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2363__B _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1758__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[11\] mod.u_arbiter.i_wb_cpu_rdt\[8\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ clknet_3_4__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2661__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1556__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[11\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1493__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2505__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2505__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2284__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2036__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1971_ _0337_ _0350_ _0366_ _0367_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2523_ mod.u_arbiter.i_wb_cpu_rdt\[22\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] _0777_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2454_ _0958_ _0745_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1405_ _0852_ _0868_ _0885_ mod.u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2385_ _0353_ _0626_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1336_ mod.u_cpu.cpu.decode.opcode\[2\] _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_mod.u_scanchain_local.scan_flop\[27\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3006_ io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1483__B1 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2684__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2338__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[59\] mod.u_scanchain_local.module_data_in\[58\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[21\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[62\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1529__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2170_ _0499_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[15\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2009__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1954_ mod.u_arbiter.i_wb_cpu_rdt\[4\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _1045_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1768__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1885_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _0288_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _0785_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ _0334_ _0341_ _0353_ _0408_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1940__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ _0308_ _0672_ _0677_ _0409_ _0679_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2299_ _0218_ _0614_ _0615_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2609__D mod.u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2248__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2133__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[26\]_D mod.u_arbiter.i_wb_cpu_rdt\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2487__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1998__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1998__B2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1670_ _1042_ _1095_ _1096_ _1097_ mod.u_arbiter.o_wb_cpu_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2175__A1 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[17\]_D mod.u_arbiter.i_wb_cpu_rdt\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2478__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2222_ _0329_ _0365_ _0543_ _0354_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2153_ mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] mod.u_arbiter.i_wb_cpu_dbus_adr\[25\]
+ _1163_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2084_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1989__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__C _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2986_ io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1937_ _0249_ _0325_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2402__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1799_ mod.u_cpu.raddr\[1\] _0227_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1913__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1591__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2469__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2840_ _2840_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__1877__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2771_ _0180_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2396__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1722_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _1127_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2745__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1653_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\]
+ _1076_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_99_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1584_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _0846_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1371__A2 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2205_ _0379_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2136_ _0481_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2067_ _0440_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2084__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2969_ io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2191__B _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2622__D _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2387__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2311__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2618__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[41\] mod.u_scanchain_local.module_data_in\[40\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[3\] clknet_3_0__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2768__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2378__A1 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__B2 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2550__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2153__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[60\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2823_ _2823_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2369__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2754_ _0163_ io_in[12] mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1705_ _1042_ _1121_ _1122_ _1123_ mod.u_arbiter.o_wb_cpu_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ _0097_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1636_ _1071_ _1067_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1567_ _0930_ _0963_ _0828_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1344__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1498_ _0837_ _0825_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2119_ mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] mod.u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _1164_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2617__D _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2057__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_126_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2141__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1583__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2296__B1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2590__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2048__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0760_ _0761_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ mod.u_cpu.rf_ram_if.rdata0\[2\] _0895_ mod.u_cpu.rf_ram_if.rtrig0 _0896_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2523__A1 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1352_ _0829_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3022_ io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1885__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2806_ _2806_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_34_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2737_ _0146_ io_in[12] mod.u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2668_ _0080_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1619_ _1053_ _1057_ _1058_ mod.u_arbiter.o_wb_cpu_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2599_ _0030_ io_in[12] mod.u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__A1 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2554__B _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1492__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _0241_ _0244_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2441__B1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1885__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ _0793_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_142_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2453_ _0863_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1404_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2384_ _0368_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1335_ _0824_ mod.u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3005_ io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1483__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1483__B2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1538__A2 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1527__C mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2338__I1 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2499__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2499__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1777__A2 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1529__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2268__C _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ _0251_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1884_ _0294_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[5\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] _0750_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2193__A2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1940__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2436_ _0259_ _0732_ _0733_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2367_ mod.u_cpu.cpu.immdec.imm30_25\[4\] _0635_ _0678_ mod.u_cpu.cpu.immdec.imm30_25\[5\]
+ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2298_ _0828_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _0218_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2651__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1931__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1695__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[17\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1922__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2279__B _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2221_ _0404_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ _0489_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2674__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2083_ _0448_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_mod.u_scanchain_local.scan_flop\[24\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2985_ io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1936_ mod.u_arbiter.i_wb_cpu_rdt\[8\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _1044_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1867_ _0280_ _0278_ _0284_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1798_ _0229_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _0247_ _0314_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1677__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[61\]_CLK clknet_3_2__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2697__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[14\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_mod.u_scanchain_local.scan_flop\[29\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ _0179_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ _1038_ _1134_ _1135_ mod.u_arbiter.o_wb_cpu_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1893__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1443__I1 mod.u_cpu.rf_ram.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1652_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _1079_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\]
+ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1583_ _0846_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_63_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1659__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2204_ _0528_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2135_ mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] mod.u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _1164_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2320__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1674__A4 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2066_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1831__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2968_ io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1919_ _0316_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2899_ _2899_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2139__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[34\] mod.u_arbiter.i_wb_cpu_rdt\[31\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2382__B _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2712__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_0__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1813__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2822_ _2822_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2369__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2753_ _0162_ io_in[12] mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1704_ mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] _1041_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2684_ _0096_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1635_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1566_ _0927_ _0964_ _0985_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2541__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1497_ _0927_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2118_ _0472_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3098_ wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ _0430_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_70_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2296__B2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2735__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2296__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2220__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ _0887_ _0018_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2523__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1351_ _0837_ _0838_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2287__B _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3021_ io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2287__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2805_ _0214_ io_in[12] mod.u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2608__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2736_ _0145_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2211__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2667_ _0079_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1618_ mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] _1042_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2598_ _0029_ io_in[12] mod.u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1549_ _0996_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2758__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[6\] mod.u_arbiter.i_wb_cpu_rdt\[3\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ clknet_3_4__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2450__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2202__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[50\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2505__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2269__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1492__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2441__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__B2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ mod.u_arbiter.i_wb_cpu_rdt\[21\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] _0777_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2452_ _0863_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0928_ _0864_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1403_ _0882_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2383_ _0249_ _0333_ _0626_ _0325_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1334_ _0824_ mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_99_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3004_ io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1483__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2719_ _0128_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1538__A3 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.input_buf_clk io_in[8] mod.u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2580__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2499__A1 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2147__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1777__A3 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ _0347_ _0348_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2414__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1883_ mod.u_arbiter.i_wb_cpu_rdt\[21\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _0288_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2504_ _0784_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2435_ _0926_ _0259_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2366_ _0669_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2297_ _0827_ _0940_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2405__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[5\]_D mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[64\] mod.u_scanchain_local.module_data_in\[63\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[26\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1729__B _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2279__C _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2220_ _0544_ _0314_ _0317_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] mod.u_arbiter.i_wb_cpu_dbus_adr\[24\]
+ _1163_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2082_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__B _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2984_ io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1935_ _0251_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1610__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1866_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _0859_ _0278_ _0283_ _0284_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1797_ _1180_ _0219_ _0227_ _0228_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2418_ _0249_ _0311_ _0719_ _0252_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2349_ _0352_ _0529_ _0627_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1365__A1 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2165__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1668__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1912__I0 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1840__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] _1038_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _1053_ _1082_ _1083_ mod.u_arbiter.o_wb_cpu_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1582_ _1023_ _1026_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1356__A1 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2203_ _0335_ _0350_ _0358_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2134_ _0480_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2791__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2065_ _0439_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2084__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1831__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2967_ io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _2898_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1918_ _0310_ _0311_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1849_ mod.u_cpu.cpu.genblk3.csr.mstatus_mpie _0261_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1347__A1 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2155__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmod.u_scanchain_local.scan_flop\[27\] mod.u_arbiter.i_wb_cpu_rdt\[24\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2664__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[14\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1510__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2066__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1813__A2 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2821_ _2821_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2752_ _0161_ io_in[12] mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1703_ _1119_ _1120_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1577__A1 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2683_ _0095_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[60\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1634_ _1067_ _1069_ _1070_ mod.u_arbiter.o_wb_cpu_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1565_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1496_ mod.u_cpu.cpu.state.o_cnt\[2\] _0928_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0947_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1371__C _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2117_ mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] mod.u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _1164_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3097_ wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2057__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2048_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\]
+ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2483__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2687__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1804__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[13\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[37\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[31\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1568__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[28\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2517__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2517__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1562__B _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2048__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2220__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1350_ mod.u_cpu.cpu.csr_d_sel _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3020_ io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1899__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2287__A2 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _0213_ io_in[12] mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2735_ _0144_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2211__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2666_ _0078_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1970__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ mod.u_cpu.cpu.o_wdata1 io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2478__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1548_ mod.u_cpu.cpu.state.o_cnt_r\[3\] _0997_ _0929_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1479_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2450__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2202__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2702__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1713__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2388__B _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2269__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[7] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2441__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2520_ _0792_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2451_ _1177_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1402_ _0858_ _0868_ _0882_ _0883_ mod.u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2382_ _0689_ _0690_ _0255_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2298__B _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1333_ mod.u_cpu.rf_ram_if.rcnt\[0\] _0822_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3003_ io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2718_ _0127_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2725__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2196__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[38\]_D mod.u_scanchain_local.module_data_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1943__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ _0062_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2499__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2163__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2423__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__A4 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2187__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2338__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _0347_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2748__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2414__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1882_ _0293_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1925__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2503_ mod.u_arbiter.i_wb_cpu_rdt\[12\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] _0750_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2434_ _0408_ _0354_ _0531_ _0341_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2365_ _0517_ _0674_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2350__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2296_ _0311_ _0570_ _0611_ _0408_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2102__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[40\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2405__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1392__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2192__I1 mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2341__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2341__B2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[57\] mod.u_scanchain_local.module_data_in\[56\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[19\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1907__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2332__B2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2332__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _0488_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_mod.u_scanchain_local.scan_flop\[63\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2081_ _0447_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2983_ io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1934_ _0327_ _0328_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2399__A1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1865_ _0952_ _0827_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1796_ mod.u_cpu.raddr\[0\] _0226_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2571__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2417_ _0315_ _0721_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2348_ _0651_ _0660_ _0661_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2279_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _0408_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2562__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2165__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2593__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2078__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] _1073_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1581_ _0830_ mod.u_cpu.cpu.bne_or_bge _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2553__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2305__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ _0333_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2133_ mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] mod.u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _1164_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1903__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_cpu.rf_ram.RAM0_CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2966_ io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2897_ _2897_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1917_ _0313_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2241__B1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1848_ _1029_ _0269_ _0270_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1779_ _1181_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2544__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__A2 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1510__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _2820_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_13_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2751_ _0160_ io_in[12] mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2682_ _0094_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1702_ _1119_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1577__A2 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] _1042_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1564_ _0987_ _0995_ _1000_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1495_ _0941_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2116_ _0471_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3096_ wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2047_ _0429_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2949_ _2949_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2214__B1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2517__A1 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2517__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1562__C _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1879__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2781__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1979__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _0212_ io_in[12] mod.u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_mod.u_scanchain_local.scan_flop\[8\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ _0143_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2665_ _0077_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1616_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _1044_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ mod.u_cpu.rf_ram_if.wdata1_r\[7\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1970__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ mod.u_cpu.cpu.decode.op26 _0841_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1478_ mod.u_cpu.cpu.state.o_cnt\[2\] _0928_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0929_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2654__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3079_ la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_126_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1961__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[6] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1952__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2450_ _0828_ _0259_ _0742_ _0743_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1401_ mod.u_cpu.cpu.immdec.imm11_7\[2\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1704__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2381_ _1046_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2677__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1332_ mod.u_cpu.rf_ram_if.rcnt\[1\] _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_mod.u_scanchain_local.scan_flop\[27\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[12\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3002_ io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[27\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__A3 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ _0126_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1943__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2648_ _0061_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2579_ _0005_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__C _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__C _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2187__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1934__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1698__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ _1181_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1622__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1881_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _0288_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2502_ _0783_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_31_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2433_ _0730_ _0534_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2364_ _0323_ _0672_ _0675_ _0251_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2350__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2295_ _0532_ _0612_ _0368_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1433__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2326__C1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2080_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2715__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2982_ io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ _0319_ _0320_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1864_ _0276_ _0278_ _0282_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1428__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1795_ mod.u_cpu.raddr\[0\] _0226_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2020__A1 mod.u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2416_ _0311_ _0334_ _0626_ _0247_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2347_ mod.u_cpu.cpu.immdec.imm30_25\[2\] _0637_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2278_ _1046_ mod.u_arbiter.i_wb_cpu_rdt\[17\] _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_77_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2562__A2 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2169__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2738__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1428__I1 mod.u_cpu.rf_ram.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2250__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1580_ _0831_ _1025_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2002__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[30\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2305__A2 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2201_ _0249_ _0251_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2132_ _0479_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2063_ _0438_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1816__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2965_ io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2896_ _2896_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2241__B2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2241__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1916_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1847_ mod.u_cpu.cpu.genblk3.csr.mie_mtie _0269_ _1036_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2529__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1778_ _1044_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2544__A2 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[53\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1991__B1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2535__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2299__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1897__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2223__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2750_ _0159_ io_in[12] mod.u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2681_ _0093_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1701_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _1108_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1632_ _1038_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1563_ _1006_ _1007_ _0205_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1494_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _0942_ _0943_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3095_ user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2115_ mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] mod.u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _1164_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1441__S mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2046_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\]
+ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2948_ _2948_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2214__B2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ _2879_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2583__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2517__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2020__B _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[32\] mod.u_arbiter.i_wb_cpu_rdt\[29\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2205__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1731__A3 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2802_ _0211_ io_in[12] mod.u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2733_ _0142_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2664_ _0076_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1615_ _1053_ _1054_ _1055_ mod.u_arbiter.o_wb_cpu_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1436__S mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2595_ mod.u_cpu.rf_ram_if.wdata1_r\[6\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1546_ mod.u_cpu.cpu.decode.op22 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1477_ mod.u_cpu.cpu.mem_bytecnt\[0\] _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2029_ _0420_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2435__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[5] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1400_ _0865_ _0846_ _0026_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_29_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2380_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[21\] _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1331_ mod.u_cpu.rf_ram_if.rcnt\[2\] _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3001_ io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2716_ _0125_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2647_ _0060_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1393__C _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2353__B1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2578_ _0004_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2621__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1529_ _0864_ _0960_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2771__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmod.u_scanchain_local.scan_flop\[4\] mod.u_arbiter.i_wb_cpu_rdt\[1\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ clknet_3_4__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[8\]_D mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__B1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1698__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_2__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _0292_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2501_ mod.u_arbiter.i_wb_cpu_rdt\[11\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] _0750_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2644__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2432_ _0245_ _0252_ _0355_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2794__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2363_ _0323_ _0310_ _0364_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2294_ _0311_ _0337_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1377__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2413__I1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2326__B1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1924__I0 mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1579__B mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1852__A2 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1604__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2667__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[11\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1368__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_mod.u_scanchain_local.scan_flop\[26\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1915__I0 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1540__A1 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2981_ io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1932_ _0310_ _0311_ _0318_ _0322_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1863_ _0278_ _0281_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1794_ _0869_ _0225_ _0226_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1359__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2020__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2159__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2415_ _0381_ _0543_ _0707_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_85_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2346_ _0408_ _0652_ _0659_ _0376_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1531__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2277_ _0251_ _0357_ _0364_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1598__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2011__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1770__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2078__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[62\] mod.u_scanchain_local.module_data_in\[61\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[24\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_1_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1589__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2002__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1761__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2200_ _0333_ _0354_ _0380_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2131_ mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] mod.u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _1164_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2062_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1816__A2 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2964_ io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1915_ mod.u_arbiter.i_wb_cpu_rdt\[6\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _1044_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ _2895_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2241__A2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2529__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1846_ _0998_ _0267_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2529__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1777_ _0843_ mod.u_cpu.cpu.state.init_done _0990_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1752__A1 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1504__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2329_ _0544_ _0529_ _0627_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1991__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__B2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1743__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2299__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A2 mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2223__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2680_ _0092_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1700_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1631_ _1065_ _1066_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1982__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1562_ mod.u_cpu.cpu.csr_d_sel _1011_ _0825_ _0926_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1734__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1493_ _0938_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ _0470_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3094_ user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2045_ _0428_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2947_ _2947_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2728__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _2878_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_50_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1973__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _0247_ _0252_ _0253_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1725__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_scanchain_local.scan_flop\[20\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A2 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2205__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[25\] mod.u_arbiter.i_wb_cpu_rdt\[22\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_142_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1964__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1964__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1731__A4 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ _0210_ io_in[12] mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ _0141_ io_in[12] mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2663_ _0075_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1944__C _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] _1042_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2594_ mod.u_cpu.rf_ram_if.wdata1_r\[5\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1545_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1516__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2380__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1476_ _0825_ _0828_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_mod.u_scanchain_local.scan_flop\[43\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3077_ la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2028_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2435__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[4] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1937__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2362__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[66\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3000_ io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2573__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__C _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1928__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2715_ _0124_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2050__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2646_ _0059_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2353__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2353__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2577_ _0003_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1528_ _0837_ _0976_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1459_ mod.u_cpu.rf_ram_if.rdata1\[6\] _0910_ _0912_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2105__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1910__S _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ mod.u_scanchain_local.clk_out io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1467__I0 mod.u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2344__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2596__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2032__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ _0782_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_10_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1494__C _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2431_ _0839_ _0390_ _0565_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2362_ _0340_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2293_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_arbiter.i_wb_cpu_rdt\[3\] _1046_ _0611_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1377__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2629_ _0042_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2326__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2326__B2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1924__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2565__A1 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1368__A2 mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2317__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__D mod.u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1931_ _0326_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ _0827_ _0933_ _0280_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0845_
+ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_35_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2761__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2556__A1 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1793_ _0221_ _0822_ _0823_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2308__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2414_ _0308_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2345_ _0408_ _0657_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1531__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1524__I mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2276_ _0357_ _0570_ _0595_ _0241_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2244__B1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1770__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2634__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[55\] mod.u_scanchain_local.module_data_in\[54\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[17\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2784__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1761__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2130_ _0478_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2061_ _0437_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2474__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2963_ io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1914_ _1181_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2894_ _2894_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2529__A1 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1845_ mod.u_cpu.cpu.decode.co_ebreak _0928_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0997_
+ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1776_ _0826_ _1176_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1455__S _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2328_ _0253_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2657__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_mod.u_scanchain_local.scan_flop\[10\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ _0315_ _0529_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_mod.u_scanchain_local.scan_flop\[25\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1440__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1339__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1630_ _1065_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1982__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1783__B _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1561_ _0830_ _1008_ _1009_ _1011_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1734__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1492_ _0926_ _0933_ mod.u_cpu.cpu.immdec.imm11_7\[0\] _0931_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1498__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2113_ mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] mod.u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _1164_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3093_ user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2044_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\]
+ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _2946_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2877_ _2877_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_31_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ mod.u_arbiter.i_wb_cpu_rdt\[1\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _1045_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1973__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1759_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[18\] mod.u_arbiter.i_wb_cpu_rdt\[15\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] clknet_3_0__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1716__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2800_ _0209_ io_in[12] mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1404__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0140_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _0074_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1613_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _1050_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2593_ mod.u_cpu.rf_ram_if.wdata1_r\[4\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1544_ _0991_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2380__A2 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1475_ mod.u_cpu.cpu.decode.opcode\[0\] _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_3__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3076_ la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2027_ _0419_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_36_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2929_ _2929_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1946__A2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[3] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2273__I mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1937__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2718__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1928__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2714_ _0123_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2645_ _0058_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[10\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2353__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2576_ _0002_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1463__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1527_ _0838_ _0976_ _0977_ mod.u_cpu.cpu.csr_d_sel _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_45_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1458_ _0917_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2105__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1389_ _0873_ mod.u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3128_ wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1467__I1 mod.u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_5__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2344__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1607__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2280__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[33\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2430_ _0837_ _0390_ _0559_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2335__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ _0310_ _0334_ _0516_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2292_ _0525_ _0608_ _0609_ _0610_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2099__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2690__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1846__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _0041_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2326__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2559_ _0814_ _1180_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1837__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[56\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2014__A1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2317__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _0327_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2253__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1861_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2005__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2556__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1792_ mod.u_cpu.rf_ram_if.rcnt\[0\] _0225_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2413_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_arbiter.i_wb_cpu_rdt\[8\] _1045_ _0719_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2308__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2344_ _0335_ _0339_ _0652_ _0252_ _0371_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2275_ _0532_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1819__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2586__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1770__A3 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2320__B _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[48\] mod.u_scanchain_local.module_data_in\[47\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[10\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2230__B _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2474__A1 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2962_ io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2226__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1913_ _1044_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2893_ _2893_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2529__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1844_ mod.u_cpu.cpu.state.o_cnt_r\[3\] mod.u_cpu.cpu.state.o_cnt\[2\] _0267_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1775_ _0827_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ _0349_ _0365_ _0623_ _0354_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1471__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2258_ _0215_ _0577_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2366__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2189_ _0514_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1440__A2 _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2601__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2456__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2751__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0830_ _1009_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1491_ _0926_ _0933_ _0931_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1498__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2112_ _0469_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3092_ la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_78_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ _0427_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2447__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2945_ _2945_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2876_ _2876_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1827_ _0249_ _0251_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1758_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2624__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1689_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] _1108_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_1_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2774__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1661__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2213__I1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2429__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[8\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0139_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _0073_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1612_ _1041_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2592_ mod.u_cpu.rf_ram_if.wdata1_r\[3\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2797__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1543_ _0929_ _0992_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[24\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1474_ _0925_ mod.u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xmod.u_scanchain_local.out_flop mod.u_scanchain_local.module_data_in\[69\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.data_out_i vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_68_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_mod.u_scanchain_local.scan_flop\[39\]_CLK clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1340__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3075_ la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2026_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _0416_ _0418_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\]
+ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1643__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2928_ _2928_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2859_ _2859_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_123_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1924__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1954__I0 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[2] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[30\] mod.u_arbiter.i_wb_cpu_rdt\[27\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] clknet_3_4__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1398__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1570__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2713_ _0122_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2050__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2644_ _0057_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2575_ _0001_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1936__I0 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1971__C _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1526_ _0975_ _0971_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1561__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1457_ mod.u_cpu.rf_ram_if.rdata1\[5\] _0907_ _0912_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1388_ mod.u_cpu.raddr\[1\] _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3127_ wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3058_ la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2009_ _0252_ _0333_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2501__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1607__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2032__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1543__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2459__I mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2291_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _0525_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2627_ _0040_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2558_ mod.u_cpu.rf_ram_if.rgnt _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2489_ mod.u_arbiter.i_wb_cpu_rdt\[6\] _0744_ _0757_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] _0750_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1509_ _0949_ _0951_ _0953_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_134_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1837__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[2\] mod.u_arbiter.i_wb_cpu_ack io_in[11] mod.u_arbiter.i_wb_cpu_dbus_sel\[0\]
+ clknet_3_0__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2014__A2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1773__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2317__A3 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1540__A4 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1860_ _0279_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2005__A2 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1791_ _1180_ _0219_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1764__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2412_ _0709_ _0713_ _0718_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2343_ _0517_ _0654_ _0656_ _0247_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2274_ _0379_ _0357_ _0527_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1819__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__B _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1469__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2244__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _0365_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1755__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[22\]_D mod.u_arbiter.i_wb_cpu_rdt\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[23\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2483__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2235__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[30\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2230__C _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2171__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[13\]_D mod.u_arbiter.i_wb_cpu_rdt\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2474__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2226__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1912_ mod.u_arbiter.i_wb_cpu_rdt\[11\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _1044_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2892_ _2892_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2405__C _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1985__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1843_ _0266_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1774_ mod.u_arbiter.i_wb_cpu_ack _1041_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1737__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[46\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2326_ _0325_ _0544_ _0336_ _0349_ _0640_ _0326_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2257_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[16\] _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2188_ _0400_ _0311_ _0332_ _0330_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1500__B mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2315__C _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1976__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1726__I _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_4__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[60\] mod.u_scanchain_local.module_data_in\[59\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[22\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1967__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2392__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[69\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1490_ _0938_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] mod.u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _1164_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3091_ la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2576__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2042_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2447__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2416__B _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2944_ _2944_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2875_ _2875_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2080__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1826_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1974__C _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1757_ _0960_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2383__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1688_ _1042_ _1108_ _1109_ _1110_ mod.u_arbiter.o_wb_cpu_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[7] mod.u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2309_ _0340_ _0515_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2438__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2374__A1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2599__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2429__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__B _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2062__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2660_ _0072_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1611_ _1049_ _1051_ _1052_ mod.u_arbiter.o_wb_cpu_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2365__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2591_ mod.u_cpu.rf_ram_if.wdata1_r\[2\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1542_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _0929_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1473_ mod.u_cpu.rf_ram_if.wdata0_r\[6\] mod.u_cpu.rf_ram_if.wdata1_r\[6\] _0865_
+ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1340__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3074_ la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_78_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2025_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2927_ _2927_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2858_ _2858_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_102_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2789_ _0198_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1809_ mod.u_cpu.cpu.genblk3.csr.timer_irq_r _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2741__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2356__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2108__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[1] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2044__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[23\] mod.u_arbiter.i_wb_cpu_rdt\[20\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1858__B1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ _0121_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2764__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2643_ _0056_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2574_ _0000_ io_in[12] mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1525_ _0975_ _0971_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1456_ _0916_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1387_ mod.u_cpu.raddr\[0\] _0870_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3126_ wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_71_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3057_ la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1616__A3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _0886_ _0345_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2026__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2329__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1552__A2 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2501__A1 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2352__I1 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2637__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2787__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[23\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2568__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2233__C _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[38\]_CLK clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1791__A2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2290_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _0218_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__B _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0039_ io_in[12] mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2557_ _1035_ _0813_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2488_ _0774_ _0775_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1508_ _0957_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1439_ _0906_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2495__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3109_ wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_93_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1773__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2325__I1 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _1035_ _0219_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1764__A2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2802__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ mod.u_cpu.cpu.immdec.imm24_20\[3\] _0714_ _0716_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ _0253_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2273_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[7] mod.u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ _0245_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2609_ mod.u_cpu.rf_ram_if.wdata0_r\[3\] io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1507__A2 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2180__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2171__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2891_ _2891_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1911_ mod.u_arbiter.i_wb_cpu_rdt\[10\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _1044_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1842_ _0261_ _0263_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1985__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1773_ _0830_ _0839_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1737__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2421__C _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2325_ mod.u_arbiter.i_wb_cpu_rdt\[26\] mod.u_arbiter.i_wb_cpu_rdt\[10\] _1045_ _0640_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2256_ mod.u_arbiter.i_wb_cpu_rdt\[0\] _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2187_ _0251_ _0332_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1673__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1425__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1976__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[1\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1361__B1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[53\] mod.u_scanchain_local.module_data_in\[52\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[15\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_95_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1967__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2392__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2110_ _0468_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3090_ la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2041_ _0426_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1655__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2943_ _2943_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1407__B2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2416__C _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2874_ _2874_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_102_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ mod.u_arbiter.i_wb_cpu_rdt\[14\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _1044_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1756_ _0826_ _0946_ _1159_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[6] mod.u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[13\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2383__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] _1041_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2308_ _0332_ _0333_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2239_ _0352_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2670__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[36\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] _1042_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2590_ mod.u_cpu.rf_ram_if.wdata1_r\[1\] io_in[12] mod.u_cpu.rf_ram_if.wdata1_r\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1541_ _0938_ mod.u_cpu.cpu.genblk3.csr.mcause31 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1472_ _0924_ mod.u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1382__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2693__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3073_ la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2024_ _1035_ _1151_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ _2926_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2857_ _2857_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1808_ _1151_ _0233_ _0234_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2788_ _0197_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2356__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1739_ _0859_ _1148_ _0990_ mod.u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1506__B _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2513__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1619__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[0] _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_scanchain_local.scan_flop\[59\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2292__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[16\] mod.u_arbiter.i_wb_cpu_rdt\[13\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_68_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1858__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0120_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2642_ _0055_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2573_ _0027_ io_in[12] mod.u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1524_ mod.u_cpu.cpu.alu.i_rs1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1455_ mod.u_cpu.rf_ram_if.rdata1\[4\] _0904_ _0912_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1386_ _0871_ mod.u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3125_ wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3056_ la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_71_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2007_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _0345_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1616__A4 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2274__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2026__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2589__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2909_ _2909_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2265__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2017__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2008__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2559__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2625_ _0038_ io_in[12] mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2556_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0944_ _0810_ _0812_ _0813_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1507_ mod.u_cpu.cpu.state.o_cnt_r\[1\] mod.u_cpu.cpu.state.o_cnt_r\[0\] mod.u_cpu.cpu.state.o_cnt_r\[3\]
+ mod.u_cpu.cpu.state.o_cnt_r\[2\] _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2487_ _1175_ _0757_ _0750_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1438_ mod.u_cpu.rf_ram.rdata\[5\] mod.u_cpu.rf_ram.data\[5\] _0026_ _0906_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__A1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3108_ wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1369_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _0824_ _0849_ mod.u_cpu.cpu.immdec.imm24_20\[2\]
+ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3039_ la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2247__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2604__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A1 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2754__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__B1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ _0308_ _0711_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2341_ _0335_ _0365_ _0623_ _0353_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_5__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ _0525_ _0590_ _0591_ _0592_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1604__B _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2477__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[6] mod.u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _0323_ _0355_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2401__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2627__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2608_ mod.u_cpu.rf_ram_if.wdata0_r\[2\] io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2539_ mod.u_arbiter.i_wb_cpu_rdt\[30\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[31\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] _0777_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2777__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1507__A3 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[22\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2468__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[1\]_D mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[37\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1691__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2300__S _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2890_ _2890_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1910_ mod.u_arbiter.i_wb_cpu_rdt\[30\] mod.u_arbiter.i_wb_cpu_rdt\[14\] _1046_ _0309_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ _0833_ _1029_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1772_ _1168_ _1172_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2324_ mod.u_cpu.cpu.immdec.imm30_25\[1\] _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1370__A1 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2255_ _0567_ _0525_ _0575_ _0576_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2186_ _0340_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1425__A2 _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1361__B2 mod.u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[46\] mod.u_scanchain_local.module_data_in\[45\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[8\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1416__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1352__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2040_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2942_ _2942_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1407__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2873_ _2873_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2080__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1824_ _1181_ mod.u_arbiter.i_wb_cpu_rdt\[15\] _0248_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1755_ _0827_ _0981_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[5] mod.u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] _1104_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1343__A1 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2307_ _0323_ _0325_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2238_ mod.u_cpu.cpu.immdec.imm19_12_20\[3\] _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1646__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] _0498_ _1163_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2115__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1954__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2531__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2531__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2062__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1540_ mod.u_cpu.cpu.decode.co_ebreak _0832_ _0988_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__1573__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ mod.u_cpu.rf_ram_if.wdata0_r\[5\] mod.u_cpu.rf_ram_if.wdata1_r\[5\] _0865_
+ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3072_ la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2925_ _2925_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2856_ _2856_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1807_ mod.u_cpu.cpu.state.ibus_cyc _0233_ _1035_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2787_ _0196_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _1141_ _1143_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1669_ mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] _1073_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2513__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2513__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2292__A2 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2044__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[9\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1858__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2283__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__B _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _0119_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2641_ _0054_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2660__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2572_ _0944_ _1035_ _1143_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1523_ _0840_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[10\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1454_ _0915_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1385_ mod.u_cpu.raddr\[0\] _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3124_ wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2006_ _0379_ _0341_ _0396_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2274__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2026__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__B _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2908_ _2908_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_143_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2839_ _2839_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__1537__A1 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[26\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2265__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2017__A2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2683__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[33\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1528__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2489__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2008__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1767__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2213__S _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2624_ _0037_ io_in[12] mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1519__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2555_ _0825_ _0827_ _1166_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[49\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2486_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _0744_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1506_ _0955_ _0956_ _0825_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1437_ _0905_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1368_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] mod.u_cpu.rf_ram_if.rtrig0 _0856_ _0857_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2495__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3107_ wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3038_ la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2123__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[25\]_D mod.u_arbiter.i_wb_cpu_rdt\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2486__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__B2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1997__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1749__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2174__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[16\]_D mod.u_arbiter.i_wb_cpu_rdt\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2340_ _0315_ _0392_ _0625_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1921__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2579__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _0525_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1988__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[5] mod.u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1986_ _0356_ _0381_ _0382_ _0244_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2401__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ mod.u_cpu.rf_ram_if.wdata0_r\[1\] io_in[12] mod.u_cpu.rf_ram_if.wdata0_r\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2538_ _0801_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2469_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _0744_ _0750_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2468__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[0\] io_in[10] io_in[11] mod.u_arbiter.o_wb_cpu_cyc
+ clknet_3_2__leaf_mod.u_scanchain_local.clk mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2721__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ mod.u_cpu.cpu.genblk3.csr.mstatus_mpie _0833_ _0262_ _0859_ _0264_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] _1173_ _1168_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2395__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ _0636_ _0638_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1370__A2 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2254_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _0376_ _0323_ _0308_ _0524_ _0576_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2185_ _0332_ _0334_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1969_ _0330_ _0349_ _0351_ _0249_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2744__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2386__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1361__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2074__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmod.u_scanchain_local.scan_flop\[39\] mod.u_scanchain_local.module_data_in\[38\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[1\] clknet_3_3__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2377__A1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2617__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2941_ _2941_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2767__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2872_ _2872_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_mod.u_scanchain_local.scan_flop\[21\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ _1044_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2368__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1754_ _0954_ mod.u_cpu.cpu.decode.opcode\[1\] _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2368__B2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[4] mod.u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[36\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _1100_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_143_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__I1 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2306_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[9\] _0408_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1343__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2237_ _0553_ _0525_ _0559_ _0560_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _0464_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2099_ _1143_ _0458_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2359__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2131__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2531__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1573__A2 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1470_ _0923_ mod.u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2125__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2022_ _0958_ _1143_ _1035_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2038__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _2924_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2855_ _2855_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1806_ _0938_ _0218_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2786_ _0195_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1737_ _0926_ _1144_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1668_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _1093_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1599_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2513__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2544__B _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1491__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1875__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0053_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2805__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ _1035_ _0821_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1522_ _0965_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1453_ mod.u_cpu.rf_ram_if.rdata1\[3\] _0901_ _0912_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1384_ _0868_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3123_ wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3054_ la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2005_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[10\] _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2274__A3 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2907_ _2907_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_143_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ _2838_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2769_ _0178_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2620__D _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1537__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1759__I _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2017__A3 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[21\] mod.u_arbiter.i_wb_cpu_rdt\[18\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2489__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2489__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ _0024_ io_in[12] mod.u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2554_ _0808_ _0811_ _1035_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1505_ _0837_ _0839_ _0831_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2485_ _0772_ _0773_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1436_ mod.u_cpu.rf_ram_if.rdata0\[5\] _0904_ mod.u_cpu.rf_ram_if.rtrig0 _0905_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1367_ mod.u_cpu.rf_ram_if.rtrig0 _0833_ _0854_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[8\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3106_ wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3037_ la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2247__A3 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[4\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1930__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1694__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[69\] mod.u_scanchain_local.module_data_in\[68\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[31\] clknet_3_3__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2650__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1921__A2 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2270_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _0218_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[4] mod.u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ _0353_ _0365_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[16\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2606_ mod.u_cpu.rf_ram_if.wtrig0 io_in[12] mod.u_cpu.rf_ram_if.genblk1.wtrig0_r
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2537_ mod.u_arbiter.i_wb_cpu_rdt\[29\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] _0777_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2468_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] _1168_ _0757_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1419_ _0894_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2399_ _0705_ _0706_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2673__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[23\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1600__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2092__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[39\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2219__I0 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0938_ _0837_ _0825_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2395__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1883__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2322_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2696__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2253_ _0256_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2184_ mod.u_cpu.cpu.immdec.imm31 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2219__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1830__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1968_ _0332_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2386__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1899_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _0288_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1433__I1 mod.u_cpu.rf_ram.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2310__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1821__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2372__B _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2940_ _2940_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2871_ _2871_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_71_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2282__B _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1822_ _0246_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2368__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1753_ mod.u_cpu.cpu.bufreg.c_r _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1684_ _1053_ _1106_ _1107_ mod.u_arbiter.o_wb_cpu_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[3] mod.u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2525__C1 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2305_ _1046_ mod.u_arbiter.i_wb_cpu_rdt\[25\] _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2236_ mod.u_cpu.cpu.immdec.imm19_12_20\[3\] _0376_ _0525_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2167_ mod.u_cpu.cpu.bufreg.i_sh_signed mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] _1143_
+ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2098_ _0960_ _1143_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2711__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2531__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[51\] mod.u_scanchain_local.module_data_in\[50\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[13\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_73_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2507__C1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3070_ la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2021_ _0886_ _0346_ _0413_ _0414_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2286__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2734__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2923_ _2923_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2854_ _2854_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2785_ _0194_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1805_ mod.u_cpu.rf_ram.regzero _0967_ _0232_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1736_ _0825_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2210__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1667_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _1093_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1598_ _1036_ mod.u_cpu.cpu.state.ibus_cyc _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2513__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2618__D _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2219_ mod.u_arbiter.i_wb_cpu_rdt\[5\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _1045_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2277__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1875__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2201__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2607__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[20\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2757__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2097__B _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[35\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1491__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ mod.u_cpu.cpu.mem_bytecnt\[1\] _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1891__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1521_ _0966_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1452_ _0914_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3122_ wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1383_ mod.u_cpu.rf_ram_if.rcnt\[0\] mod.u_cpu.rf_ram_if.rcnt\[1\] mod.u_cpu.rf_ram_if.rcnt\[2\]
+ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3053_ la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2259__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2004_ _1045_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _2906_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2431__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2837_ _2837_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2768_ _0177_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2699_ _0108_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1719_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2137__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2364__C _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[14\] mod.u_arbiter.i_wb_cpu_rdt\[11\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2489__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2489__A1 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2622_ _0023_ io_in[12] mod.u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2553_ _0926_ _0809_ _0810_ _0827_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1504_ _0828_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2484_ mod.u_arbiter.i_wb_cpu_rdt\[4\] _0744_ _0750_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1435_ _0887_ _0021_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2449__C _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1366_ mod.u_cpu.cpu.decode.op26 mod.u_cpu.cpu.decode.co_ebreak _0829_ _0840_ _0855_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3105_ wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3036_ la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2404__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[4\]_D mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1694__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2375__B _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2269__C _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[3] mod.u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2398__B1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1984_ _0379_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2605_ _0035_ io_in[12] mod.u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2536_ _0800_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_103_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2467_ _1168_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1418_ mod.u_cpu.rf_ram.rdata\[1\] mod.u_cpu.rf_ram.data\[1\] _0026_ _0894_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2398_ mod.u_cpu.cpu.immdec.imm24_20\[3\] _0686_ _0687_ mod.u_cpu.cpu.immdec.imm24_20\[2\]
+ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1676__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1349_ mod.u_cpu.cpu.bne_or_bge _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2389__B1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1667__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_cpu.rf_ram.RAM0_CEN _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1911__I0 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2092__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2325__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[7\]_CLK clknet_3_1__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1355__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2321_ _0258_ _0634_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _0351_ _0568_ _0570_ _0349_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2155__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1658__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2183_ _0510_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _0249_ _0325_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2386__A3 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1594__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1898_ _0301_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2519_ mod.u_arbiter.i_wb_cpu_rdt\[20\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] _0777_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2640__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1346__A1 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2790__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2074__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2145__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1821__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1958__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ _2870_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_15_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ _0242_ _0243_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2663__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ mod.u_cpu.cpu.alu.i_rs1 _1155_ _1156_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1683_ mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] _1073_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[2] mod.u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[13\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2525__B1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2525__C2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2304_ _0990_ _0619_ _0620_ _0374_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2235_ _0390_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2166_ _0496_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1500__A1 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ mod.u_cpu.cpu.state.o_cnt_r\[1\] mod.u_cpu.cpu.state.o_cnt_r\[0\] _0929_ _0458_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2473__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2300__I0 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2999_ io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[29\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1552__B _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__I _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2383__B _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[44\] mod.u_scanchain_local.module_data_in\[43\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[6\] clknet_3_4__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2686__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[36\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1558__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_7__f_mod.u_scanchain_local.clk_I clknet_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2507__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1730__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _0259_ _0346_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1889__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2922_ _2922_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2853_ _2853_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2784_ _0193_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ mod.u_cpu.rf_ram.regzero _0824_ _0232_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1735_ _0954_ mod.u_arbiter.i_wb_cpu_dbus_we _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2210__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1666_ _1042_ _1092_ _1093_ _1094_ mod.u_arbiter.o_wb_cpu_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1564__A4 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1597_ _1040_ mod.u_arbiter.o_wb_cpu_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2468__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ _0528_ _0529_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2277__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2149_ mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] mod.u_arbiter.i_wb_cpu_dbus_adr\[23\]
+ _1163_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1788__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2201__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1520_ _0933_ _0968_ _0969_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1451_ mod.u_cpu.rf_ram_if.rdata1\[2\] _0898_ _0912_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2701__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1382_ _0868_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3121_ wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3052_ la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2003_ _0883_ _0390_ _0345_ _0397_ _0398_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2905_ _2905_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2431__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2836_ _2836_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2767_ _0176_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2698_ _0107_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1718_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _1127_
+ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_mod.u_scanchain_local.scan_flop\[37\]_D mod.u_scanchain_local.module_data_in\[36\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1649_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _1079_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1942__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2198__B _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2422__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2153__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2724__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2186__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[28\]_D mod.u_arbiter.i_wb_cpu_rdt\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2489__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2621_ _0022_ io_in[12] mod.u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ _0944_ _1143_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1503_ _0926_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2483_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _1168_ _0757_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1434_ _0903_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1365_ mod.u_cpu.cpu.immdec.imm24_20\[1\] _0847_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3104_ wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3035_ la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2101__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2747__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2819_ _2819_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[34\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1391__A2 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[49\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2340__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1906__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__C _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1897__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[2] mod.u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2398__A1 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1983_ _0323_ _0251_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2604_ _0034_ io_in[12] mod.u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2535_ mod.u_arbiter.i_wb_cpu_rdt\[28\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] _0777_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2570__A1 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2466_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] mod.u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1417_ _0892_ _0893_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2322__A1 mod.u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2397_ _0308_ _0699_ _0704_ _0409_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_mod.u_scanchain_local.scan_flop\[62\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1348_ _0830_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3018_ io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2086__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2389__B2 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2561__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2552__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2320_ mod.u_cpu.cpu.immdec.imm30_25\[1\] _0390_ _0632_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1355__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2251_ _0337_ _0350_ _0571_ _0572_ _0368_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2304__B2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2304__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2182_ mod.u_cpu.cpu.genblk3.csr.timer_irq_r _0236_ _0238_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2592__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2068__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1966_ _0253_ _0244_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1594__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1897_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0288_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2518_ _0791_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2449_ _0341_ _0381_ _0395_ _0376_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2161__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_6__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0241_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1751_ mod.u_cpu.cpu.alu.i_rs1 mod.u_cpu.cpu.bufreg.c_r _1155_ _1156_ _1157_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1682_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] _1104_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[1] mod.u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2525__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2303_ _0940_ _0990_ _0376_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1923__B _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2234_ _0408_ _0333_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2165_ mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] mod.u_arbiter.i_wb_cpu_dbus_adr\[31\]
+ _1163_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1887__I0 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1500__A2 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2096_ _0452_ _0457_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2998_ io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1949_ _1044_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[6\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2383__C _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[37\] mod.u_scanchain_local.module_data_in\[36\]
+ io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1558__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2507__A1 mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1494__A1 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2921_ _2921_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2443__B1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2630__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1797__A2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2852_ _2852_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2783_ _0192_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1803_ _0024_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2780__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1734_ _0825_ _0827_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1665_ mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] _1073_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1596_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _1038_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ mod.u_cpu.cpu.immdec.imm19_12_20\[1\] _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2277__A3 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2148_ _0487_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1485__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2079_ _0446_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[7\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1960__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1712__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1476__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2653__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2394__B _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1738__B _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1400__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1951__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ _0913_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1381_ _0866_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2288__C _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3120_ wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3051_ la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2002_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _0345_ _0218_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2904_ _2904_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _2835_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_91_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_mod.u_scanchain_local.scan_flop\[19\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2766_ _0175_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2697_ _0106_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1717_ _1053_ _1131_ _1132_ mod.u_arbiter.o_wb_cpu_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1648_ _1053_ _1079_ _1080_ _1081_ mod.u_arbiter.o_wb_cpu_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1942__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1579_ _0837_ _1025_ mod.u_cpu.cpu.bne_or_bge _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2676__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[26\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[9\] mod.u_arbiter.i_wb_cpu_rdt\[6\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ clknet_3_1__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1558__B mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1933__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2408__I mod.u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ _0021_ io_in[12] mod.u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2551_ _0838_ _0508_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2699__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2482_ _1168_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1502_ _0843_ mod.u_cpu.cpu.state.init_done _0952_ _0828_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1433_ mod.u_cpu.rf_ram.rdata\[4\] mod.u_cpu.rf_ram.data\[4\] _0026_ _0903_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1688__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1364_ _0850_ _0851_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1423__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3103_ wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3034_ la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2818_ _2818_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2749_ _0158_ io_in[12] mod.u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2002__B _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2340__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1851__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2095__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[1] mod.u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _0325_ _0329_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ _0033_ io_in[12] mod.u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2534_ _0799_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1418__S _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2465_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1416_ mod.u_cpu.rf_ram_if.rdata0\[1\] _0824_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2396_ _0371_ _0701_ _0702_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2322__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1347_ mod.u_cpu.cpu.decode.co_ebreak _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3017_ io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2714__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1833__A1 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2010__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1364__A3 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2159__S _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[67\] mod.u_scanchain_local.module_data_in\[66\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[29\] clknet_3_2__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1824__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2001__B2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2001__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2552__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1355__A3 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _0544_ _0543_ _0513_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _0990_ _0508_ _0509_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2737__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1815__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[33\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1965_ _0339_ _0350_ _0362_ _0244_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1418__I1 mod.u_cpu.rf_ram.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[48\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2240__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1896_ _0300_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xmod.u_scanchain_local.output_buffers\[2\] mod.u_scanchain_local.data_out_i mod.u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__2240__B2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2517_ mod.u_arbiter.i_wb_cpu_rdt\[19\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] _0777_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_2448_ _0408_ _0314_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2379_ _0540_ _0688_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1806__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2231__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2519__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2298__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2352__S _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1750_ _0827_ _0954_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2222__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[52\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2222__B2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1681_ _1042_ _1103_ _1104_ _1105_ mod.u_arbiter.o_wb_cpu_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_mod.u_cpu.rf_ram.RAM0_A[0] mod.u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2525__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2302_ mod.u_cpu.cpu.immdec.imm7 _0390_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2289__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2233_ _0247_ _0251_ _0341_ _0556_ _0408_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2164_ _0495_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2095_ _0455_ _0456_ _0436_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1431__S mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1948_ _0218_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1879_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _0288_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2010__B _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2452__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2582__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2507__A2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2920_ _2920_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2443__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2443__B2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2851_ _2851_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2782_ _0191_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1802_ _0231_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1733_ _0957_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1664_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\]
+ _1085_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1595_ _1039_ mod.u_arbiter.o_wb_cpu_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1426__S mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2216_ _0521_ _0525_ _0540_ _0541_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2147_ mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] mod.u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _1163_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1485__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2078_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2434__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2434__B2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1960__A3 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1476__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A1 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1738__C _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1400__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ mod.u_cpu.rf_ram_if.rcnt\[0\] _0822_ _0823_ mod.u_cpu.rf_ram_if.wen0_r _0867_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3050_ la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2001_ _0255_ _0394_ _0396_ _0357_ _0376_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2416__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _2903_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2834_ _2834_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2765_ _0174_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1716_ mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] _1073_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2696_ _0105_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_mod.u_scanchain_local.scan_flop\[5\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1647_ mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] _1073_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1578_ mod.u_cpu.cpu.csr_d_sel _0975_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_mod.u_scanchain_local.scan_flop\[7\]_D mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2620__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2770__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2550_ _0944_ mod.u_cpu.cpu.ctrl.i_jump _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _1170_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1501_ mod.u_cpu.cpu.genblk3.csr.o_new_irq _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1432_ _0902_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1363_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _0824_ _0849_ mod.u_cpu.cpu.immdec.imm24_20\[3\]
+ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3102_ wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3033_ la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1503__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2817_ _2817_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_30_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2748_ _0157_ io_in[12] mod.u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2643__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2679_ _0091_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2793__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[12\] mod.u_arbiter.i_wb_cpu_rdt\[9\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ clknet_3_5__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1367__A1 mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2095__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_cpu.rf_ram.RAM0_D[0] mod.u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _0346_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2666__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2602_ mod.u_cpu.rf_ram_if.rtrig0 io_in[12] mod.u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2533_ mod.u_arbiter.i_wb_cpu_rdt\[27\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] _0777_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2464_ _0753_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1415_ _0887_ mod.u_cpu.rf_ram_if.rtrig0 _0017_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2395_ _0341_ _0626_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1346_ mod.u_cpu.cpu.decode.op21 _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1530__A1 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3016_ io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2086__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1833__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2010__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2239__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1824__A2 mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1588__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2537__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2537__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ mod.u_cpu.cpu.alu.cmp_r _0990_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1815__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _0249_ _0351_ _0361_ _0252_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1579__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1895_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0288_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2516_ _0790_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1751__A1 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2447_ _0933_ _0390_ _0741_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2378_ mod.u_cpu.cpu.immdec.imm24_20\[1\] _0686_ _0687_ mod.u_cpu.cpu.immdec.imm24_20\[0\]
+ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1806__A2 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1847__B _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2519__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2519__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1990__B2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2298__A2 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2222__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] _1041_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1981__A1 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2704__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2301_ _0618_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2232_ _0512_ _0554_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2163_ mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] mod.u_arbiter.i_wb_cpu_dbus_adr\[30\]
+ _1163_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _0454_ _0930_ _0986_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2461__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1947_ _0990_ _1147_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1878_ _0291_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1724__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2452__A2 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2727__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1963__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[32\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[47\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2443__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2850_ _2850_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1801_ _1036_ mod.u_cpu.rf_ram_if.rreq_r _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2781_ _0190_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1732_ mod.u_cpu.cpu.state.init_done mod.u_cpu.cpu.genblk3.csr.o_new_irq _1142_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1663_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] _1088_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1594_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2215_ mod.u_cpu.cpu.immdec.imm19_12_20\[1\] _0259_ _0525_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2146_ _0486_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ _0445_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2434__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1397__B _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2979_ io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2198__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1945__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[42\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1476__A3 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[42\] mod.u_scanchain_local.module_data_in\[41\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[4\] clknet_3_0__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_77_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1400__A3 _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2361__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2000_ _0254_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2902_ _2902_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2416__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2833_ _2833_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2764_ _0173_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1715_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1927__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2695_ _0104_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] _1076_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1577_ mod.u_cpu.cpu.csr_d_sel mod.u_cpu.cpu.csr_imm _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[65\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2104__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2129_ mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] mod.u_arbiter.i_wb_cpu_dbus_adr\[13\]
+ _1164_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2407__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1918__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2040__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1394__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2343__B2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2343__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1765__B _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1909__A1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2480_ _0768_ _0769_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1500_ mod.u_cpu.cpu.csr_d_sel mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] mod.u_cpu.cpu.state.init_done
+ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1431_ mod.u_cpu.rf_ram_if.rdata0\[4\] _0901_ mod.u_cpu.rf_ram_if.rtrig0 _0902_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2334__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2334__B2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3101_ wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1362_ mod.u_cpu.rf_ram_if.rtrig0 _0848_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2595__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3032_ la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2816_ _2816_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_20_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ _0156_ io_in[12] mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2678_ _0090_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1629_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _1056_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2564__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1367__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2316__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[4\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ mod.u_cpu.cpu.immdec.imm11_7\[2\] _0376_ _0308_ _0335_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2601_ _0032_ io_in[12] mod.u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2532_ _0798_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2555__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1358__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2463_ _0577_ _0744_ _0750_ _0751_ _0755_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2307__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1414_ _0891_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2394_ _0245_ _0693_ _0352_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1345_ mod.u_cpu.cpu.decode.op26 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1530__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3015_ io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2610__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2546__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2760__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2537__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1334__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2633__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ _0321_ _0355_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1894_ _0299_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2783__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2515_ mod.u_arbiter.i_wb_cpu_rdt\[18\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] _0777_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2446_ _0368_ _0721_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2377_ _0258_ _0685_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2216__B1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2519__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2656__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1430__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1981__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2300_ _0617_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _0525_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2231_ _0353_ _0543_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2162_ _0494_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2093_ mod.u_cpu.cpu.ctrl.i_jump _0964_ _0453_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2995_ io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1946_ _0307_ _0344_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ mod.u_arbiter.i_wb_cpu_rdt\[18\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _0288_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1972__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1724__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2679__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1903__S _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2429_ _0838_ _0390_ _0551_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1488__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__B1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1412__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1963__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1479__A1 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1612__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1651__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0225_ _0230_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2780_ _0189_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ _0874_ _0878_ _0883_ _0886_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1662_ _1053_ _1090_ _1091_ mod.u_arbiter.o_wb_cpu_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1593_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2214_ _0533_ _0538_ _0539_ _0308_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2145_ mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] mod.u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _1163_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2076_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\]
+ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2978_ io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1929_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1945__A2 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[35\] mod.u_scanchain_local.module_data_in\[34\]
+ io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] clknet_3_1__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2361__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2901_ _2901_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ _2832_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2763_ _0172_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1714_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _1127_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1927__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2694_ _0014_ io_in[12] mod.u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] _1076_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ _0987_ _0995_ _1000_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1453__S _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2104__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2717__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2128_ _0477_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2059_ _0417_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1615__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[31\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1918__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[46\]_CLK clknet_3_5__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1909__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1337__I _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ _0887_ _0020_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1361_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _0824_ _0849_ mod.u_cpu.cpu.immdec.imm24_20\[4\]
+ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2334__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2098__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3031_ la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1845__A1 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2270__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2815_ _2815_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[32\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2746_ _0155_ io_in[12] mod.u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2677_ _0089_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1628_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1559_ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _0863_
+ _0864_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1911__S _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1836__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[7\] mod.u_arbiter.i_wb_cpu_rdt\[4\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ clknet_3_1__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1827__A1 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_mod.u_scanchain_local.scan_flop\[55\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2252__B2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2451__I _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2004__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _0031_ io_in[12] mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2531_ mod.u_arbiter.i_wb_cpu_rdt\[26\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] _0777_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2555__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2462_ _0751_ _1168_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2307__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1413_ _0888_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2393_ _0252_ _0699_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1344_ mod.u_cpu.cpu.decode.op21 _0829_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3014_ io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1818__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__A1 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2729_ _0138_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2482__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2234__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2585__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2537__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1899__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__D mod.u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1350__I mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _0349_ _0355_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2225__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ mod.u_arbiter.i_wb_cpu_rdt\[26\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0288_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2514_ _0789_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2445_ _0247_ _0249_ _0408_ _0313_ _0258_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2376_ _0218_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1461__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2519__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[3\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[65\] mod.u_scanchain_local.module_data_in\[64\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[27\] clknet_3_3__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2455__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2207__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__B _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1430__A2 _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _0314_ _0400_ _0311_ _0330_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2600__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] mod.u_arbiter.i_wb_cpu_dbus_adr\[29\]
+ _1163_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2092_ _0859_ _0833_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2446__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2750__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2994_ io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1945_ _0308_ _0309_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1876_ _0290_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2428_ _0540_ _0729_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ _1046_ mod.u_arbiter.i_wb_cpu_rdt\[29\] _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1488__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2437__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__B2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2623__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2773__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1479__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_opt_1_1_mod.u_scanchain_local.clk clknet_opt_1_0_mod.u_scanchain_local.clk
+ clknet_opt_1_1_mod.u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__B1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1730_ _0863_ _1140_ _0837_ mod.u_arbiter.i_wb_cpu_dbus_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1661_ mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] _1073_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1592_ _1036_ mod.u_cpu.cpu.state.ibus_cyc _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2213_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_arbiter.i_wb_cpu_rdt\[4\] _1046_ _0539_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2144_ _0485_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2075_ _0444_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2419__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2977_ io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2646__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1928_ _1045_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_mod.u_scanchain_local.scan_flop\[7\]_SI mod.u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1859_ _0277_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1633__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmod.u_scanchain_local.scan_flop\[28\] mod.u_arbiter.i_wb_cpu_rdt\[25\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] clknet_3_4__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1397__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2212__C _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2900_ _2900_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2669__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2831_ _2831_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_2762_ _0171_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1713_ _1053_ _1128_ _1129_ mod.u_arbiter.o_wb_cpu_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2693_ _0103_ io_in[12] mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1644_ _1053_ _1076_ _1077_ _1078_ mod.u_arbiter.o_wb_cpu_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_99_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ _1022_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1560__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] mod.u_arbiter.i_wb_cpu_dbus_adr\[12\]
+ _1164_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2058_ _0435_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2040__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.output_buffers\[3\]_I clknet_opt_1_1_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2223__B _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1790__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1360_ _0824_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2596__D mod.u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2098__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3030_ la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2270__A2 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2814_ _2814_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_20_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2022__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2745_ _0154_ io_in[12] mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ _0088_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1627_ _1053_ _1063_ _1064_ mod.u_arbiter.o_wb_cpu_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1558_ _0838_ _0928_ mod.u_cpu.cpu.mem_bytecnt\[1\] _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1533__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1489_ mod.u_cpu.cpu.immdec.imm31 _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1772__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1827__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2707__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1348__I _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _0797_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2461_ _0752_ _1168_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1763__A1 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1412_ _0889_ _0866_ _0867_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2392_ _0323_ _0315_ _0562_ _0380_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[30\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1343_ mod.u_cpu.cpu.csr_d_sel _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3013_ io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_mod.u_scanchain_local.scan_flop\[30\]_D mod.u_arbiter.i_wb_cpu_rdt\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_mod.u_scanchain_local.scan_flop\[45\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1818__A2 mod.u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1459__S _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2243__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ _0137_ io_in[12] mod.u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2659_ _0071_ io_in[12] mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2234__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1993__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[10\] mod.u_arbiter.i_wb_cpu_rdt\[7\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ clknet_3_4__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_52_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[12\]_D mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[22\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2473__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ _0356_ _0350_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _0298_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1984__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ mod.u_arbiter.i_wb_cpu_rdt\[17\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] _0750_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1736__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2444_ _0738_ _0739_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2375_ _0829_ _1145_ _0958_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2216__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1975__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1727__A1 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[45\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[58\] mod.u_scanchain_local.module_data_in\[57\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[20\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1966__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2160_ _0493_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2091_ mod.u_cpu.cpu.ctrl.i_jump _1006_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2993_ io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1944_ _0331_ _0338_ _0342_ _0258_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1875_ mod.u_arbiter.i_wb_cpu_rdt\[17\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _0288_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1709__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[68\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ mod.u_cpu.cpu.decode.co_ebreak _0259_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ _0256_ _0668_ _0670_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1488__A3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2289_ _0310_ _0570_ _0604_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2575__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2437__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2316__B _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2070__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1948__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1559__S0 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1939__B2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] _1088_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1591_ _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2364__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2598__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2212_ _0535_ _0536_ _0537_ _0364_ _0256_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2143_ mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] mod.u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _1163_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2074_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2419__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[2\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2976_ io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2052__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1927_ _0323_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1467__S _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1858_ _0938_ _0846_ _0929_ _0991_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2355__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ _1180_ _0224_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1469__I0 mod.u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2346__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ _2830_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_56_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2034__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2761_ _0170_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1712_ mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] _1073_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2692_ _0102_ io_in[12] mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1643_ mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] _1073_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1574_ mod.u_cpu.rf_ram.rdata\[7\] mod.u_cpu.rf_ram.data\[7\] _0026_ _1022_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2126_ _0476_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2057_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] _0434_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2959_ io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2763__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1379__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2328__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1551__A2 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[40\] mod.u_scanchain_local.module_data_in\[39\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[2\] clknet_3_0__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_142_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2567__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__A1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1790__A2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1542__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2636__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2465__I _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__A3 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2786__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ _2813_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0153_ io_in[12] mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ _0087_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1626_ mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] _1042_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1781__A2 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1557_ mod.u_cpu.cpu.mem_if.signbit _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1488_ _0825_ _0827_ mod.u_cpu.cpu.csr_d_sel _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] mod.u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _1164_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3089_ la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_74_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__A3 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2659__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2237__B1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_2__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2460_ _0949_ _0747_ _1177_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1763__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1411_ mod.u_cpu.rf_ram.data\[0\] _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2391_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_arbiter.i_wb_cpu_rdt\[6\] _1045_ _0699_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1515__A2 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1342_ _0830_ mod.u_cpu.cpu.bne_or_bge _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3012_ io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2228__B1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _0136_ io_in[12] mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2658_ _0070_ io_in[12] mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2801__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1609_ _1038_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2589_ mod.u_cpu.cpu.o_wen0 io_in[12] mod.u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1681__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1960_ _0310_ _0311_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1891_ mod.u_arbiter.i_wb_cpu_rdt\[25\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _0288_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _0788_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_143_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2443_ _0825_ _0259_ _0308_ _0352_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2374_ _0344_ _0683_ _0684_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1727__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1966__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_mod.u_scanchain_local.scan_flop\[44\]_CLK clknet_3_4__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[0\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_mod.u_scanchain_local.scan_flop\[59\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] _0416_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2992_ io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1943_ _0332_ _0340_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1957__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1874_ _0289_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2426_ _0697_ _0728_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2357_ mod.u_cpu.cpu.immdec.imm30_25\[3\] _0637_ _0665_ _0308_ _0669_ mod.u_cpu.cpu.immdec.imm30_25\[4\]
+ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_85_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2288_ _0325_ _0371_ _0606_ _0218_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1948__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[12\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2373__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1559__S1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1462__I _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ io_in[9] _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2364__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2211_ _0354_ _0365_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2521__C1 mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2142_ _0484_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2073_ _0443_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1627__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2975_ io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[35\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[14\] _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1857_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _0276_ _0845_ _0277_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2355__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1788_ _0219_ _0223_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2409_ _0715_ _0686_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1469__I1 mod.u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2346__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__A1 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1609__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_mod.u_scanchain_local.scan_flop\[58\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2760_ _0169_ io_in[12] mod.u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1711_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2691_ _0016_ io_in[12] mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1642_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _1067_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\]
+ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2337__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1573_ _0865_ _1020_ _1021_ mod.u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1848__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2125_ mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] mod.u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _1164_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ _0415_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2958_ io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1909_ _0258_ _0255_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2889_ _2889_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_68_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2264__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[33\] mod.u_arbiter.i_wb_cpu_rdt\[30\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2588__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2016__A1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2319__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[1\]_CLK clknet_3_3__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__A4 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2812_ _2812_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_108_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2007__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2743_ _0152_ io_in[12] mod.u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0086_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1625_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _1060_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2430__B _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1556_ _0828_ _0954_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1487_ mod.u_cpu.cpu.bufreg2.i_cnt_done _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2108_ _1139_ _0460_ _0467_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3088_ la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2039_ _0425_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_51_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2246__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2730__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1936__S _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1763__A3 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ _0866_ _0867_ mod.u_cpu.rf_ram.rdata\[0\] _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2603__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2390_ _0697_ _0698_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1341_ mod.u_cpu.cpu.decode.co_mem_word _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3011_ io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2753__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2726_ _0135_ io_in[12] mod.u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2657_ _0013_ io_in[12] mod.u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1608_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1046_
+ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2588_ mod.u_cpu.cpu.o_wen1 io_in[12] mod.u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1539_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2467__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[0\]_D io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmod.u_scanchain_local.scan_flop\[5\] mod.u_arbiter.i_wb_cpu_rdt\[2\] io_in[11] mod.u_arbiter.i_wb_cpu_dbus_sel\[3\]
+ clknet_3_4__leaf_mod.u_scanchain_local.clk mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2335__B _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__B1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2776__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1890_ _0297_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2511_ mod.u_arbiter.i_wb_cpu_rdt\[16\] _0778_ _0756_ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] _0750_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2442_ _0390_ _0255_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2373_ mod.u_cpu.cpu.immdec.imm30_25\[5\] _0637_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2449__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1672__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2649__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2709_ _0118_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2799__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1360__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1415__A2 mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_1_1_mod.u_scanchain_local.clk_I clknet_opt_1_0_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1351__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1654__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1942_ _0253_ _0247_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1873_ mod.u_arbiter.i_wb_cpu_rdt\[16\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1957__A3 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2425_ mod.u_cpu.cpu.decode.op21 _0259_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1342__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2356_ _0218_ _0634_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2287_ _0215_ mod.u_arbiter.i_wb_cpu_rdt\[2\] _0407_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1956__I0 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1581__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmod.u_scanchain_local.scan_flop\[63\] mod.u_scanchain_local.module_data_in\[62\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[25\] clknet_3_6__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1572__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2210_ _0354_ _0527_ _0241_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2141_ mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] mod.u_arbiter.i_wb_cpu_dbus_adr\[19\]
+ _1163_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2521__C2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2072_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] _0434_ _0436_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2974_ io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1925_ _1044_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2052__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1856_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1787_ _0220_ _0222_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1991__C _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1563__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2408_ mod.u_cpu.cpu.immdec.imm24_20\[4\] _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2339_ _0353_ _0529_ _0627_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__A2 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1618__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[43\]_CLK clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2291__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[58\]_CLK clknet_3_6__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1554__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2503__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2503__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2034__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1710_ _1124_ _1119_ _1120_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2690_ _0015_ io_in[12] mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1641_ _1075_ _1071_ _1065_ _1066_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_67_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1572_ _0865_ mod.u_cpu.rf_ram_if.wdata1_r\[7\] _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2124_ _0475_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2055_ _0433_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_74_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1986__C _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2957_ io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2888_ _2888_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1908_ mod.u_cpu.cpu.bufreg.i_sh_signed _0259_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1839_ _0996_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2016__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[26\] mod.u_arbiter.i_wb_cpu_rdt\[23\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] clknet_3_5__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1775__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1527__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[25\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_mod.u_scanchain_local.clk clknet_0_mod.u_scanchain_local.clk clknet_3_7__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2255__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ _2811_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2007__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2742_ _0151_ io_in[12] mod.u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1766__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ _0085_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1624_ _1059_ _1061_ _1062_ mod.u_arbiter.o_wb_cpu_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1555_ _1004_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.scan_flop\[33\]_D mod.u_arbiter.i_wb_cpu_rdt\[30\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1486_ mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2107_ _0460_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3087_ la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2038_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2246__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2113__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1509__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_mod.u_scanchain_local.scan_flop\[48\]_SE io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[24\]_D mod.u_arbiter.i_wb_cpu_rdt\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2237__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1996__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1748__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1340_ _0826_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2173__A1 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_mod.u_scanchain_local.scan_flop\[15\]_D mod.u_arbiter.i_wb_cpu_rdt\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3010_ io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2492__I _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2228__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1987__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1739__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0134_ io_in[12] mod.u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2656_ _0069_ io_in[12] mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1607_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1046_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2587_ _0028_ io_in[12] mod.u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1538_ mod.u_cpu.cpu.state.o_cnt_r\[1\] mod.u_cpu.cpu.state.o_cnt_r\[0\] mod.u_cpu.cpu.state.o_cnt_r\[3\]
+ mod.u_cpu.cpu.state.o_cnt_r\[2\] _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2578__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1469_ mod.u_cpu.rf_ram_if.wdata0_r\[4\] mod.u_cpu.rf_ram_if.wdata1_r\[4\] _0865_
+ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1571__I _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[0\]_CLK clknet_3_2__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1969__B2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1969__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2510_ _0787_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2394__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ _0244_ _0251_ _0736_ _0381_ _0368_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2720__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2372_ mod.u_cpu.cpu.immdec.imm7 _1156_ _0669_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2449__A2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2082__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2708_ _0117_ io_in[12] mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2602__D mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2385__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0052_ io_in[12] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1515__B _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2376__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1351__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_mod.u_scanchain_local.out_flop_D mod.u_scanchain_local.module_data_in\[69\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2151__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2990_ io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2064__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ _0333_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1872_ _0216_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1957__A4 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1386__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2424_ _0997_ _0390_ _0705_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2355_ _0517_ _0664_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1342__A2 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2286_ _1046_ mod.u_arbiter.i_wb_cpu_rdt\[18\] _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2616__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2766__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2358__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2121__S _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1581__A2 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmod.u_scanchain_local.scan_flop\[56\] mod.u_scanchain_local.module_data_in\[55\]
+ io_in[11] mod.u_arbiter.o_wb_cpu_adr\[18\] clknet_3_7__leaf_mod.u_scanchain_local.clk
+ mod.u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2046__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2349__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1572__A2 mod.u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__A1 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2639__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0483_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2071_ _0442_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_35_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2789__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1883__I0 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2973_ io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1924_ mod.u_arbiter.i_wb_cpu_rdt\[15\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _1045_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1855_ _0275_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1786_ _0221_ mod.u_cpu.rf_ram_if.rcnt\[1\] _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2407_ _0376_ _0685_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2338_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_arbiter.i_wb_cpu_rdt\[11\] _1045_ _0652_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2269_ _0408_ _0579_ _0589_ _0258_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2028__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1955__S _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2503__A1 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__B1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1640_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1571_ _1020_ mod.u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2123_ mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] mod.u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _1164_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _0416_ _0418_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1481__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2956_ io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2887_ _2887_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1907_ _1035_ _0306_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1838_ _0833_ _0999_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2804__CLK io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1769_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2610__D mod.u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1536__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2497__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__C2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2421__B1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmod.u_scanchain_local.scan_flop\[19\] mod.u_arbiter.i_wb_cpu_rdt\[16\] io_in[11]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] clknet_3_0__leaf_mod.u_scanchain_local.clk
+ mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1775__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2810_ _2810_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2741_ _0150_ io_in[12] mod.u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1766__A2 mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ _0084_ io_in[12] mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1623_ mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] _1042_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_mod.u_scanchain_local.scan_flop\[42\]_CLK clknet_3_0__leaf_mod.u_scanchain_local.clk
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1554_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r _1005_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1485_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

