// This is the unpowered netlist.
module serv_0 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_arbiter.o_wb_cpu_adr[0] ;
 wire \u_arbiter.o_wb_cpu_adr[10] ;
 wire \u_arbiter.o_wb_cpu_adr[11] ;
 wire \u_arbiter.o_wb_cpu_adr[12] ;
 wire \u_arbiter.o_wb_cpu_adr[13] ;
 wire \u_arbiter.o_wb_cpu_adr[14] ;
 wire \u_arbiter.o_wb_cpu_adr[15] ;
 wire \u_arbiter.o_wb_cpu_adr[16] ;
 wire \u_arbiter.o_wb_cpu_adr[17] ;
 wire \u_arbiter.o_wb_cpu_adr[18] ;
 wire \u_arbiter.o_wb_cpu_adr[19] ;
 wire \u_arbiter.o_wb_cpu_adr[1] ;
 wire \u_arbiter.o_wb_cpu_adr[20] ;
 wire \u_arbiter.o_wb_cpu_adr[21] ;
 wire \u_arbiter.o_wb_cpu_adr[22] ;
 wire \u_arbiter.o_wb_cpu_adr[23] ;
 wire \u_arbiter.o_wb_cpu_adr[24] ;
 wire \u_arbiter.o_wb_cpu_adr[25] ;
 wire \u_arbiter.o_wb_cpu_adr[26] ;
 wire \u_arbiter.o_wb_cpu_adr[27] ;
 wire \u_arbiter.o_wb_cpu_adr[28] ;
 wire \u_arbiter.o_wb_cpu_adr[29] ;
 wire \u_arbiter.o_wb_cpu_adr[2] ;
 wire \u_arbiter.o_wb_cpu_adr[30] ;
 wire \u_arbiter.o_wb_cpu_adr[31] ;
 wire \u_arbiter.o_wb_cpu_adr[3] ;
 wire \u_arbiter.o_wb_cpu_adr[4] ;
 wire \u_arbiter.o_wb_cpu_adr[5] ;
 wire \u_arbiter.o_wb_cpu_adr[6] ;
 wire \u_arbiter.o_wb_cpu_adr[7] ;
 wire \u_arbiter.o_wb_cpu_adr[8] ;
 wire \u_arbiter.o_wb_cpu_adr[9] ;
 wire \u_arbiter.o_wb_cpu_cyc ;
 wire \u_arbiter.o_wb_cpu_we ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.addr[0] ;
 wire \u_cpu.rf_ram.addr[1] ;
 wire \u_cpu.rf_ram.addr[2] ;
 wire \u_cpu.rf_ram.addr[3] ;
 wire \u_cpu.rf_ram.addr[4] ;
 wire \u_cpu.rf_ram.addr[5] ;
 wire \u_cpu.rf_ram.addr[6] ;
 wire \u_cpu.rf_ram.addr[7] ;
 wire \u_cpu.rf_ram.data[0] ;
 wire \u_cpu.rf_ram.data[1] ;
 wire \u_cpu.rf_ram.data[2] ;
 wire \u_cpu.rf_ram.data[3] ;
 wire \u_cpu.rf_ram.data[4] ;
 wire \u_cpu.rf_ram.data[5] ;
 wire \u_cpu.rf_ram.data[6] ;
 wire \u_cpu.rf_ram.data[7] ;
 wire \u_cpu.rf_ram.i_wdata[0] ;
 wire \u_cpu.rf_ram.i_wdata[1] ;
 wire \u_cpu.rf_ram.i_wdata[2] ;
 wire \u_cpu.rf_ram.i_wdata[3] ;
 wire \u_cpu.rf_ram.i_wdata[4] ;
 wire \u_cpu.rf_ram.i_wdata[5] ;
 wire \u_cpu.rf_ram.i_wdata[6] ;
 wire \u_cpu.rf_ram.i_wdata[7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.clk ;
 wire \u_scanchain_local.clk_out ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.data_out_i ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1539_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1540_ (.I(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1541_ (.I(\u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1542_ (.A1(_1020_),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1543_ (.I(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1544_ (.I(_1024_),
    .Z(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1545_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1546_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1547_ (.A1(_1025_),
    .A2(_1026_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1548_ (.I(_1023_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1549_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1550_ (.I(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1551_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1552_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1553_ (.I(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1554_ (.I(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1555_ (.A1(_1030_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1556_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1557_ (.A1(_1035_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1558_ (.I(_1036_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1559_ (.A1(_1029_),
    .A2(\u_cpu.cpu.decode.op21 ),
    .A3(_1034_),
    .A4(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1560_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1561_ (.I(\u_cpu.cpu.decode.op21 ),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1562_ (.A1(_1040_),
    .A2(\u_cpu.cpu.decode.op26 ),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1563_ (.A1(_1029_),
    .A2(_1037_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1564_ (.A1(_1034_),
    .A2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1565_ (.A1(_1039_),
    .A2(_1041_),
    .B(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1566_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1567_ (.I(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1568_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1569_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1570_ (.A1(_1048_),
    .A2(_1031_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1571_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_1049_),
    .A3(_1042_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1572_ (.A1(_1047_),
    .A2(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1573_ (.A1(_1046_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1574_ (.A1(_1044_),
    .A2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1575_ (.A1(_1038_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1576_ (.A1(_1023_),
    .A2(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1577_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_1027_),
    .B1(_1055_),
    .B2(\u_cpu.cpu.immdec.imm24_20[3] ),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1578_ (.I(_1024_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1579_ (.A1(_1057_),
    .A2(_1054_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1580_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_1027_),
    .B1(_1055_),
    .B2(\u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1581_ (.A1(_1056_),
    .A2(_1058_),
    .A3(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1582_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_1053_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1583_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_1034_),
    .A4(_1042_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1584_ (.A1(_1024_),
    .A2(_1038_),
    .A3(_1061_),
    .A4(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1585_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_1057_),
    .B(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1586_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_1027_),
    .B1(_1055_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1587_ (.A1(_1047_),
    .A2(_1045_),
    .A3(_1050_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1588_ (.A1(_1041_),
    .A2(_1044_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1589_ (.A1(_1066_),
    .A2(_1067_),
    .B(_1023_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1590_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_1023_),
    .B1(_1055_),
    .B2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .C(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1591_ (.A1(_1064_),
    .A2(_1065_),
    .A3(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1592_ (.A1(_1060_),
    .A2(_1070_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1593_ (.I(_1027_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1594_ (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1595_ (.I(net2),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1596_ (.A1(_1072_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1597_ (.I(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1598_ (.I(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1599_ (.A1(_1071_),
    .A2(_1075_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1600_ (.I(_1076_),
    .Z(\u_arbiter.o_wb_cpu_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1601_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_1073_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1602_ (.I(_1077_),
    .Z(\u_arbiter.o_wb_cpu_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1603_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1604_ (.I(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1605_ (.I(_1079_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1606_ (.I(_1080_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1607_ (.I(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1608_ (.I(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1609_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1610_ (.A1(_1083_),
    .A2(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1611_ (.A1(_1083_),
    .A2(_1084_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1612_ (.A1(_1075_),
    .A2(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1613_ (.A1(_1072_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1614_ (.I(_1088_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1615_ (.I(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1616_ (.I(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1617_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1618_ (.A1(_1085_),
    .A2(_1087_),
    .B(_1092_),
    .ZN(\u_arbiter.o_wb_cpu_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1619_ (.I(_1089_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1620_ (.I(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1621_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_1086_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1622_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .A2(_1091_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1623_ (.A1(_1094_),
    .A2(_1095_),
    .B(_1096_),
    .ZN(\u_arbiter.o_wb_cpu_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1624_ (.A1(_1083_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(_1084_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1625_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1626_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .A2(_1091_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1627_ (.A1(_1094_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(\u_arbiter.o_wb_cpu_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1628_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _1629_ (.A1(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1630_ (.A1(_1100_),
    .A2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1631_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .A2(_1091_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1632_ (.A1(_1094_),
    .A2(_1102_),
    .B(_1103_),
    .ZN(\u_arbiter.o_wb_cpu_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1633_ (.A1(_1100_),
    .A2(_1101_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1634_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_1100_),
    .A3(_1101_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1635_ (.A1(_1075_),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1636_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .A2(_1091_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1637_ (.A1(_1104_),
    .A2(_1106_),
    .B(_1107_),
    .ZN(\u_arbiter.o_wb_cpu_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1638_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_1105_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1639_ (.I(_1090_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1640_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1641_ (.A1(_1094_),
    .A2(_1108_),
    .B(_1110_),
    .ZN(\u_arbiter.o_wb_cpu_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1642_ (.I(_1090_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1643_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1644_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_1101_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1645_ (.A1(_1112_),
    .A2(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1646_ (.A1(_1112_),
    .A2(_1113_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1647_ (.I(_1089_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1648_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .A2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1649_ (.A1(_1111_),
    .A2(_1114_),
    .A3(_1115_),
    .B(_1117_),
    .ZN(\u_arbiter.o_wb_cpu_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1650_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_1115_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1651_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1652_ (.A1(_1119_),
    .A2(_1112_),
    .A3(_1113_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1653_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .A2(_1116_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1654_ (.A1(_1111_),
    .A2(_1118_),
    .A3(_1120_),
    .B(_1121_),
    .ZN(\u_arbiter.o_wb_cpu_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1655_ (.I(_1090_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1656_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .A2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1657_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1658_ (.A1(_1124_),
    .A2(_1120_),
    .B(_1093_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1659_ (.A1(_1124_),
    .A2(_1120_),
    .B(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1660_ (.A1(_1123_),
    .A2(_1126_),
    .ZN(\u_arbiter.o_wb_cpu_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1661_ (.A1(_1124_),
    .A2(_1120_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1662_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1663_ (.A1(_1119_),
    .A2(_1112_),
    .A3(_1113_),
    .A4(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1664_ (.I(_1089_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1665_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1666_ (.A1(_1111_),
    .A2(_1127_),
    .A3(_1129_),
    .B(_1131_),
    .ZN(\u_arbiter.o_wb_cpu_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1667_ (.I(_1093_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1668_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1669_ (.A1(_1133_),
    .A2(_1129_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1670_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_1109_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1671_ (.A1(_1132_),
    .A2(_1134_),
    .B(_1135_),
    .ZN(\u_arbiter.o_wb_cpu_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1672_ (.A1(_1133_),
    .A2(_1129_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1673_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_1133_),
    .A3(_1129_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1674_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_1130_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1675_ (.A1(_1111_),
    .A2(_1136_),
    .A3(_1137_),
    .B(_1138_),
    .ZN(\u_arbiter.o_wb_cpu_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1676_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .A2(_1122_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1677_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1678_ (.A1(_1140_),
    .A2(_1137_),
    .B(_1093_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1679_ (.A1(_1140_),
    .A2(_1137_),
    .B(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1680_ (.A1(_1139_),
    .A2(_1142_),
    .ZN(\u_arbiter.o_wb_cpu_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1681_ (.A1(_1140_),
    .A2(_1137_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1682_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1683_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_1129_),
    .A4(_1144_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1684_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .A2(_1130_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1685_ (.A1(_1122_),
    .A2(_1143_),
    .A3(_1145_),
    .B(_1146_),
    .ZN(\u_arbiter.o_wb_cpu_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1686_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1687_ (.A1(_1147_),
    .A2(_1145_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1688_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(_1148_),
    .S(_1074_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1689_ (.I(_1149_),
    .Z(\u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1690_ (.A1(_1147_),
    .A2(_1145_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1691_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_1147_),
    .A3(_1145_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1692_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_1130_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1693_ (.A1(_1122_),
    .A2(_1150_),
    .A3(_1151_),
    .B(_1152_),
    .ZN(\u_arbiter.o_wb_cpu_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1694_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_1151_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1695_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(_1153_),
    .S(_1074_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1696_ (.I(_1154_),
    .Z(\u_arbiter.o_wb_cpu_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1697_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1698_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A4(_1145_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1699_ (.A1(_1155_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1700_ (.A1(_1155_),
    .A2(_1156_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1701_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_1130_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1702_ (.A1(_1122_),
    .A2(_1157_),
    .A3(_1158_),
    .B(_1159_),
    .ZN(\u_arbiter.o_wb_cpu_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1703_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1704_ (.A1(_1160_),
    .A2(_1157_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1705_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .A2(_1109_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1706_ (.A1(_1132_),
    .A2(_1161_),
    .B(_1162_),
    .ZN(\u_arbiter.o_wb_cpu_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1707_ (.A1(_1160_),
    .A2(_1157_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1708_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1709_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .A2(_1109_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1710_ (.A1(_1132_),
    .A2(_1164_),
    .B(_1165_),
    .ZN(\u_arbiter.o_wb_cpu_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1711_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_1160_),
    .A3(_1157_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1712_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1713_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .A2(_1109_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1714_ (.A1(_1132_),
    .A2(_1167_),
    .B(_1168_),
    .ZN(\u_arbiter.o_wb_cpu_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1715_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1716_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A4(_1157_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1717_ (.A1(_1169_),
    .A2(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1718_ (.I(_1090_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1719_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1720_ (.A1(_1132_),
    .A2(_1171_),
    .B(_1173_),
    .ZN(\u_arbiter.o_wb_cpu_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1721_ (.I(_1093_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_1169_),
    .A2(_1170_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1723_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1724_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_1172_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1725_ (.A1(_1174_),
    .A2(_1176_),
    .B(_1177_),
    .ZN(\u_arbiter.o_wb_cpu_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1726_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_1169_),
    .A3(_1170_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1727_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1728_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_1172_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1729_ (.A1(_1174_),
    .A2(_1179_),
    .B(_1180_),
    .ZN(\u_arbiter.o_wb_cpu_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1730_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1731_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A4(_1170_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1732_ (.A1(_1181_),
    .A2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1733_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .A2(_1172_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1734_ (.A1(_1174_),
    .A2(_1183_),
    .B(_1184_),
    .ZN(\u_arbiter.o_wb_cpu_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1735_ (.A1(_1181_),
    .A2(_1182_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1736_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1737_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_1172_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1738_ (.A1(_1174_),
    .A2(_1186_),
    .B(_1187_),
    .ZN(\u_arbiter.o_wb_cpu_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1739_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_1181_),
    .A3(_1182_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1740_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1741_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_1116_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1742_ (.A1(_1174_),
    .A2(_1189_),
    .B(_1190_),
    .ZN(\u_arbiter.o_wb_cpu_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1743_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A4(_1182_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1744_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1745_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_1116_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1746_ (.A1(_1111_),
    .A2(_1192_),
    .B(_1193_),
    .ZN(\u_arbiter.o_wb_cpu_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1747_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_1191_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1748_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A3(_1191_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1749_ (.A1(_1074_),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_1116_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1751_ (.A1(_1194_),
    .A2(_1196_),
    .B(_1197_),
    .ZN(\u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1752_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_1195_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1753_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A2(_1074_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1754_ (.A1(_1075_),
    .A2(_1198_),
    .B(_1199_),
    .ZN(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1755_ (.A1(\u_cpu.rf_ram_if.wen1_r ),
    .A2(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1756_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_1021_),
    .A3(_1022_),
    .A4(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1757_ (.A1(_1200_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1758_ (.I(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1759_ (.I(_1203_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1760_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1761_ (.A1(_1204_),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1762_ (.A1(_1032_),
    .A2(_1037_),
    .A3(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1763_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1764_ (.A1(_1207_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1765_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1766_ (.A1(\u_cpu.rf_ram.data[0] ),
    .A2(_1200_),
    .A3(_1201_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1767_ (.I(_1200_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1768_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_1021_),
    .A3(_1022_),
    .A4(\u_cpu.rf_ram_if.wen0_r ),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1769_ (.A1(_1211_),
    .A2(_1212_),
    .B(\u_cpu.rf_ram.rdata[0] ),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1770_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1771_ (.A1(_1210_),
    .A2(_1213_),
    .B(\u_cpu.rf_ram.regzero ),
    .C(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1772_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(_1214_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1773_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1774_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1775_ (.A1(\u_cpu.cpu.decode.opcode[2] ),
    .A2(\u_cpu.cpu.decode.opcode[0] ),
    .A3(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1776_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1218_),
    .A3(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1777_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_1219_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1778_ (.A1(\u_cpu.cpu.decode.opcode[2] ),
    .A2(_1031_),
    .A3(\u_cpu.cpu.csr_d_sel ),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1779_ (.A1(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1780_ (.A1(_1217_),
    .A2(_1220_),
    .A3(_1221_),
    .B(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1781_ (.A1(_1204_),
    .A2(_1224_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1782_ (.A1(_1209_),
    .A2(_1215_),
    .A3(_1216_),
    .B(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1783_ (.A1(_1206_),
    .A2(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(_1207_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1785_ (.A1(_1208_),
    .A2(_1227_),
    .B(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1786_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1787_ (.I(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1788_ (.I(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1789_ (.I0(_1206_),
    .I1(_1229_),
    .S(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1790_ (.I(_1233_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1791_ (.I(_1066_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1792_ (.I(\u_cpu.cpu.bne_or_bge ),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1793_ (.I(_1035_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1794_ (.I(_1028_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1795_ (.I(_1207_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1796_ (.I(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1797_ (.A1(_1237_),
    .A2(\u_cpu.cpu.csr_imm ),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1798_ (.A1(_1237_),
    .A2(_1239_),
    .B(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1799_ (.A1(_1236_),
    .A2(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1800_ (.A1(_1215_),
    .A2(_1216_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1801_ (.I(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1802_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1803_ (.I(\u_cpu.cpu.mem_bytecnt[1] ),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1804_ (.A1(_1246_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1805_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_1043_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1806_ (.A1(_1244_),
    .A2(_1245_),
    .A3(_1247_),
    .A4(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1807_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1808_ (.A1(_1217_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1809_ (.A1(_1250_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1810_ (.A1(_1040_),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_1043_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1811_ (.A1(_1231_),
    .A2(_1253_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1812_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .A2(_1250_),
    .B(_1252_),
    .C(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1813_ (.I(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1814_ (.A1(_1044_),
    .A2(_1243_),
    .B1(_1249_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1815_ (.I(_1035_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1816_ (.A1(_1258_),
    .A2(_1235_),
    .B(_1241_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1817_ (.A1(_1235_),
    .A2(_1242_),
    .B1(_1257_),
    .B2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(_1234_),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1819_ (.I(_1052_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1820_ (.A1(_1071_),
    .A2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1821_ (.A1(_1261_),
    .A2(_1263_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1822_ (.I(_1031_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1823_ (.I(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1824_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1825_ (.I(_1025_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1826_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.init_done ),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1827_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A3(_1031_),
    .A4(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1828_ (.A1(\u_cpu.cpu.decode.co_mem_word ),
    .A2(_1028_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1829_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1830_ (.A1(\u_cpu.cpu.branch_op ),
    .A2(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1831_ (.A1(_1036_),
    .A2(_1270_),
    .A3(_1272_),
    .B(_1048_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1832_ (.A1(_1230_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1833_ (.A1(_1269_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1834_ (.A1(_1035_),
    .A2(_1030_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1835_ (.A1(_1028_),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .B(_1276_),
    .C(\u_cpu.cpu.state.init_done ),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1836_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1837_ (.A1(_1275_),
    .A2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1838_ (.A1(_1267_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1839_ (.I(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1840_ (.A1(_1281_),
    .A2(_1247_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1841_ (.A1(_1264_),
    .A2(\u_arbiter.i_wb_cpu_dbus_we ),
    .B1(_1039_),
    .B2(_1049_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1842_ (.A1(_1271_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1843_ (.A1(_1219_),
    .A2(_1283_),
    .A3(_1284_),
    .B(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1844_ (.I(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1845_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1286_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _1846_ (.A1(_1269_),
    .A2(_1274_),
    .B1(_1277_),
    .B2(\u_cpu.cpu.state.stage_two_req ),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1847_ (.A1(_1025_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1848_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1849_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_1290_),
    .B(_1224_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1850_ (.A1(_1048_),
    .A2(_1271_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1851_ (.A1(_1264_),
    .A2(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1852_ (.I0(_1289_),
    .I1(_1291_),
    .S(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1853_ (.A1(_1287_),
    .A2(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1854_ (.A1(_1282_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1855_ (.A1(_1265_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1856_ (.A1(_1266_),
    .A2(_1280_),
    .B(_1297_),
    .C(_1052_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1857_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1858_ (.A1(_1299_),
    .A2(_1206_),
    .A3(_1226_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1859_ (.A1(_1042_),
    .A2(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1860_ (.I(_1226_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1861_ (.A1(_1258_),
    .A2(_1239_),
    .A3(_1302_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1862_ (.A1(_1239_),
    .A2(_1302_),
    .B(\u_cpu.cpu.bne_or_bge ),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1863_ (.A1(_1239_),
    .A2(_1302_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1864_ (.A1(_1237_),
    .A2(_1303_),
    .A3(_1304_),
    .A4(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1865_ (.A1(_1281_),
    .A2(_1247_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1866_ (.A1(_1258_),
    .A2(_1029_),
    .A3(\u_cpu.cpu.alu.cmp_r ),
    .A4(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1867_ (.A1(_1289_),
    .A2(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1868_ (.I(_1030_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1869_ (.A1(_1310_),
    .A2(_1272_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1870_ (.A1(_1301_),
    .A2(_1306_),
    .A3(_1309_),
    .B(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1871_ (.A1(_1293_),
    .A2(_1282_),
    .A3(_1295_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1872_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1873_ (.I(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1874_ (.A1(_1236_),
    .A2(_1246_),
    .B1(_1315_),
    .B2(_1037_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1875_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1876_ (.I0(_1317_),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(\u_cpu.cpu.bufreg.lsb[0] ),
    .S1(_1026_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1877_ (.A1(_1316_),
    .A2(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1878_ (.A1(_1314_),
    .A2(_1316_),
    .B(_1319_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1879_ (.I(_1048_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1880_ (.I(_1271_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1881_ (.A1(_1237_),
    .A2(_1319_),
    .B(_1320_),
    .C(_1321_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1882_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1883_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1884_ (.A1(_1323_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_1250_),
    .C(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1885_ (.A1(_1071_),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1886_ (.A1(_1325_),
    .A2(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1887_ (.A1(_1265_),
    .A2(_1321_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1888_ (.A1(_1327_),
    .A2(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1889_ (.A1(_0041_),
    .A2(_1322_),
    .B(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1890_ (.A1(_1257_),
    .A2(_1312_),
    .A3(_1313_),
    .A4(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1891_ (.A1(_1066_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1892_ (.A1(_1298_),
    .A2(_1332_),
    .ZN(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1893_ (.A1(_1210_),
    .A2(_1213_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1894_ (.I(_1203_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1895_ (.I0(\u_cpu.rf_ram.rdata[1] ),
    .I1(\u_cpu.rf_ram.data[1] ),
    .S(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1896_ (.I(_1334_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1897_ (.I0(\u_cpu.rf_ram.rdata[2] ),
    .I1(\u_cpu.rf_ram.data[2] ),
    .S(_1333_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1898_ (.I(_1335_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1899_ (.I0(\u_cpu.rf_ram.rdata[3] ),
    .I1(\u_cpu.rf_ram.data[3] ),
    .S(_1333_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1900_ (.I(_1336_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1901_ (.I0(\u_cpu.rf_ram.rdata[4] ),
    .I1(\u_cpu.rf_ram.data[4] ),
    .S(_1333_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1902_ (.I(_1337_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1903_ (.I0(\u_cpu.rf_ram.rdata[5] ),
    .I1(\u_cpu.rf_ram.data[5] ),
    .S(_1333_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1904_ (.I(_1338_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1905_ (.I0(\u_cpu.rf_ram.rdata[6] ),
    .I1(\u_cpu.rf_ram.data[6] ),
    .S(_1203_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1906_ (.I(_1339_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1907_ (.I0(\u_cpu.rf_ram.rdata[7] ),
    .I1(\u_cpu.rf_ram.data[7] ),
    .S(net8),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1908_ (.I(_1340_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1909_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1910_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1911_ (.I0(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .S(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1912_ (.I(_1343_),
    .Z(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1913_ (.I0(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .S(_1342_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1914_ (.I(_1344_),
    .Z(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1915_ (.I0(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .S(_1342_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1916_ (.I(_1345_),
    .Z(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1917_ (.I0(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .S(_1342_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1918_ (.I(_1346_),
    .Z(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1919_ (.I0(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .S(_1342_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1920_ (.I(_1347_),
    .Z(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1921_ (.I0(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .S(_1341_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1922_ (.I(_1348_),
    .Z(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1923_ (.I0(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .S(_1341_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1924_ (.I(_1349_),
    .Z(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _1925_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1926_ (.I0(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .I1(\u_cpu.cpu.o_wdata0 ),
    .S(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1927_ (.I(_1351_),
    .Z(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1928_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1929_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1930_ (.A1(_1353_),
    .A2(_0018_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1931_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1932_ (.I0(\u_cpu.rf_ram_if.rdata1[1] ),
    .I1(_1354_),
    .S(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1933_ (.I(_1356_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1934_ (.A1(_1353_),
    .A2(_0019_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1935_ (.I0(\u_cpu.rf_ram_if.rdata1[2] ),
    .I1(_1357_),
    .S(_1355_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1936_ (.I(_1358_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1937_ (.A1(_1353_),
    .A2(_0020_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1938_ (.I0(\u_cpu.rf_ram_if.rdata1[3] ),
    .I1(_1359_),
    .S(_1355_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1939_ (.I(_1360_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1940_ (.A1(_1353_),
    .A2(_0021_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1941_ (.I0(\u_cpu.rf_ram_if.rdata1[4] ),
    .I1(_1361_),
    .S(_1355_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1942_ (.I(_1362_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1943_ (.A1(_1352_),
    .A2(_0022_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1944_ (.I0(\u_cpu.rf_ram_if.rdata1[5] ),
    .I1(_1363_),
    .S(_1355_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1945_ (.I(_1364_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1946_ (.A1(_1352_),
    .A2(_0023_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1947_ (.I0(\u_cpu.rf_ram_if.rdata1[6] ),
    .I1(_1365_),
    .S(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1948_ (.I(_1366_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1949_ (.A1(_1210_),
    .A2(_1213_),
    .B(\u_cpu.rf_ram.regzero ),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1950_ (.I0(\u_cpu.rf_ram_if.rdata0[1] ),
    .I1(_1367_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1951_ (.I(_1368_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1952_ (.I0(\u_cpu.rf_ram_if.rdata0[2] ),
    .I1(_1354_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1953_ (.I(_1369_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1954_ (.I0(\u_cpu.rf_ram_if.rdata0[3] ),
    .I1(_1357_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1955_ (.I(_1370_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1956_ (.I0(\u_cpu.rf_ram_if.rdata0[4] ),
    .I1(_1359_),
    .S(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1957_ (.I(_1371_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1958_ (.I0(\u_cpu.rf_ram_if.rdata0[5] ),
    .I1(_1361_),
    .S(_1057_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1959_ (.I(_1372_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1960_ (.I0(\u_cpu.rf_ram_if.rdata0[6] ),
    .I1(_1363_),
    .S(_1057_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1961_ (.I(_1373_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1962_ (.I0(\u_cpu.rf_ram_if.rdata0[7] ),
    .I1(_1365_),
    .S(_1057_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1963_ (.I(_1374_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1964_ (.A1(_1020_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1965_ (.A1(_1202_),
    .A2(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1966_ (.A1(\u_cpu.raddr[0] ),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1967_ (.I(_1377_),
    .Z(\u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1968_ (.A1(\u_cpu.raddr[0] ),
    .A2(_1376_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1969_ (.A1(\u_cpu.raddr[1] ),
    .A2(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1970_ (.I(_1379_),
    .Z(\u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _1971_ (.I(_1202_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1972_ (.A1(_1041_),
    .A2(_1234_),
    .B(_1350_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1973_ (.A1(\u_cpu.cpu.immdec.imm11_7[0] ),
    .A2(_1341_),
    .A3(_1262_),
    .B(_1380_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _1974_ (.A1(_1069_),
    .A2(_1380_),
    .B1(_1381_),
    .B2(_1382_),
    .ZN(\u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1975_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_1341_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1976_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_1350_),
    .B(net8),
    .C(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1977_ (.A1(_1064_),
    .A2(net8),
    .B1(_1384_),
    .B2(_1234_),
    .ZN(\u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1978_ (.A1(_1350_),
    .A2(_1066_),
    .A3(_1202_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1979_ (.I(\u_cpu.cpu.immdec.imm11_7[2] ),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _1980_ (.A1(_1065_),
    .A2(_1380_),
    .B1(_1385_),
    .B2(_1386_),
    .ZN(\u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1981_ (.I(_1385_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1982_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1983_ (.A1(_1056_),
    .A2(_1380_),
    .B(_1388_),
    .ZN(\u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1984_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _1985_ (.A1(_1059_),
    .A2(_1380_),
    .B1(_1385_),
    .B2(_1389_),
    .ZN(\u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1986_ (.A1(_1058_),
    .A2(net8),
    .B(_1387_),
    .ZN(\u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1987_ (.I(_1236_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1988_ (.I(_1026_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1989_ (.A1(_0215_),
    .A2(_0216_),
    .B1(_1037_),
    .B2(_1267_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1990_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(_1281_),
    .A3(_1244_),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1991_ (.I(_0218_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1992_ (.A1(_1320_),
    .A2(_1266_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1993_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_0219_),
    .A3(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1994_ (.A1(_0217_),
    .A2(_0221_),
    .B(_1094_),
    .ZN(\u_arbiter.o_wb_cpu_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1995_ (.A1(_1209_),
    .A2(_1075_),
    .ZN(\u_arbiter.o_wb_cpu_we ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1996_ (.I(\u_cpu.cpu.decode.opcode[1] ),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1997_ (.A1(_1264_),
    .A2(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1998_ (.I(_1271_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1999_ (.A1(_1264_),
    .A2(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2000_ (.A1(_1207_),
    .A2(\u_cpu.cpu.bufreg.c_r ),
    .A3(_0223_),
    .A4(_0225_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2001_ (.A1(_1207_),
    .A2(_0223_),
    .A3(_0225_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2002_ (.A1(\u_cpu.cpu.bufreg.c_r ),
    .A2(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2003_ (.A1(_1321_),
    .A2(_0222_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2004_ (.A1(_0229_),
    .A2(_1284_),
    .B(_1307_),
    .C(_1265_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2005_ (.A1(_1310_),
    .A2(_1224_),
    .A3(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2006_ (.A1(_0228_),
    .A2(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2007_ (.I(_1279_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2008_ (.A1(_0226_),
    .A2(_0232_),
    .B(_0233_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2009_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1286_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2010_ (.A1(_1293_),
    .A2(_1291_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2011_ (.A1(_1293_),
    .A2(_1280_),
    .B(_0235_),
    .C(_1287_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2012_ (.A1(_1268_),
    .A2(_1273_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2013_ (.A1(_1231_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2014_ (.A1(_0234_),
    .A2(_0236_),
    .B(_0238_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2015_ (.A1(_1071_),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2016_ (.A1(_1325_),
    .A2(_1326_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2017_ (.A1(_0239_),
    .A2(_0240_),
    .B(_0238_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2018_ (.A1(_1053_),
    .A2(_0219_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2019_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A3(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2020_ (.A1(_1321_),
    .A2(_1204_),
    .B(_1328_),
    .C(_1310_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2021_ (.I(_0237_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2022_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_0241_),
    .B(_0242_),
    .C(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2023_ (.A1(_1234_),
    .A2(_0244_),
    .B(_0219_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2024_ (.A1(_1235_),
    .A2(_1025_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2025_ (.A1(_1026_),
    .A2(_0245_),
    .B(_0215_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2026_ (.A1(_1025_),
    .A2(_0216_),
    .B(_0215_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2027_ (.A1(_0216_),
    .A2(_0245_),
    .B(_0215_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2028_ (.I(net2),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2029_ (.I(_0246_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2030_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2031_ (.I(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2032_ (.I(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2033_ (.I(_0250_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2034_ (.A1(net12),
    .A2(_1073_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2035_ (.A1(_0251_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_0252_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2036_ (.I(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2037_ (.A1(_1045_),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_0254_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2038_ (.A1(_0247_),
    .A2(_0255_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2039_ (.A1(_1236_),
    .A2(_1048_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2040_ (.A1(_1268_),
    .A2(_1273_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2041_ (.A1(_0256_),
    .A2(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2042_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A4(net39),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2043_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2044_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2045_ (.A1(_1217_),
    .A2(_1276_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2046_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_0262_),
    .B(_0258_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2047_ (.A1(_0258_),
    .A2(_0261_),
    .B(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2048_ (.A1(_1258_),
    .A2(_1029_),
    .A3(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2049_ (.A1(net12),
    .A2(_1088_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2050_ (.I(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2051_ (.A1(_1310_),
    .A2(_0265_),
    .B(_0267_),
    .C(_1033_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2052_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_1046_),
    .A3(_0218_),
    .A4(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2053_ (.A1(_0255_),
    .A2(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2054_ (.A1(_1020_),
    .A2(_0270_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2055_ (.I(_1020_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2056_ (.A1(_0271_),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2057_ (.A1(_1375_),
    .A2(_0270_),
    .A3(_0272_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2058_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2059_ (.A1(\u_cpu.raddr[0] ),
    .A2(_0272_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2060_ (.A1(_0255_),
    .A2(_0269_),
    .A3(_0273_),
    .A4(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2061_ (.I(_0275_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2062_ (.A1(\u_cpu.raddr[1] ),
    .A2(_0273_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2063_ (.A1(_0270_),
    .A2(_0276_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2064_ (.I(_1217_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2065_ (.A1(_0277_),
    .A2(_0257_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2066_ (.A1(_0246_),
    .A2(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2067_ (.I(_0279_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2068_ (.A1(_1244_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2069_ (.A1(_1244_),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2070_ (.A1(_0246_),
    .A2(_0280_),
    .A3(_0281_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2071_ (.I(_1072_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2072_ (.A1(_1315_),
    .A2(_0281_),
    .B(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2073_ (.A1(_1315_),
    .A2(_0281_),
    .B(_0283_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2074_ (.A1(_1315_),
    .A2(_0281_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2075_ (.A1(_1246_),
    .A2(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2076_ (.A1(_0247_),
    .A2(_0285_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2077_ (.A1(net2),
    .A2(_1217_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2078_ (.I(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2079_ (.A1(_1244_),
    .A2(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2080_ (.I(\u_cpu.rf_ram_if.rgnt ),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2081_ (.A1(_0289_),
    .A2(_0269_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2082_ (.A1(_0282_),
    .A2(_0219_),
    .A3(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2083_ (.A1(_0288_),
    .A2(_0291_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2084_ (.A1(_0282_),
    .A2(_1281_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2085_ (.I(_0292_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2086_ (.A1(_0247_),
    .A2(_1323_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2087_ (.A1(_1072_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2088_ (.I(_0293_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2089_ (.A1(_1045_),
    .A2(_0287_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2090_ (.A1(_0217_),
    .A2(_0220_),
    .A3(_0032_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2091_ (.A1(_0294_),
    .A2(_0295_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2092_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_0287_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2093_ (.I(_1321_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2094_ (.A1(_1258_),
    .A2(_1237_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2095_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_1028_),
    .B(_1035_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2096_ (.A1(_1238_),
    .A2(_1226_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2097_ (.A1(_1239_),
    .A2(_1302_),
    .B(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2098_ (.A1(_1229_),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2099_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_1307_),
    .B(_1300_),
    .C(_0298_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2100_ (.A1(_0298_),
    .A2(_0302_),
    .B(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2101_ (.A1(_1235_),
    .A2(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2102_ (.A1(_0297_),
    .A2(_0305_),
    .B(_0032_),
    .C(_1266_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2103_ (.A1(_0296_),
    .A2(_0306_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2104_ (.A1(_1246_),
    .A2(_1290_),
    .A3(_0039_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2105_ (.I(_0307_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2106_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_0287_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2107_ (.A1(_0247_),
    .A2(_0278_),
    .B(_0308_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2108_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B(\u_cpu.cpu.mem_bytecnt[0] ),
    .C(\u_cpu.cpu.bufreg.lsb[0] ),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2110_ (.A1(_1231_),
    .A2(_0309_),
    .A3(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2111_ (.A1(_0256_),
    .A2(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2112_ (.I(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2113_ (.I(_0258_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2114_ (.A1(_1317_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2115_ (.A1(_0313_),
    .A2(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2116_ (.I(_0258_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2117_ (.I(_0266_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2118_ (.A1(net39),
    .A2(_0317_),
    .B(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2119_ (.A1(net12),
    .A2(_1089_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2120_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2121_ (.A1(_0320_),
    .A2(_0313_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2122_ (.I(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2123_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_0321_),
    .B1(_0323_),
    .B2(_1317_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2124_ (.A1(_0316_),
    .A2(_0319_),
    .B(_0324_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2125_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_0314_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2126_ (.A1(_1317_),
    .A2(net39),
    .B(_0314_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2127_ (.A1(_0313_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2128_ (.A1(net39),
    .A2(_0316_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2129_ (.A1(_0325_),
    .A2(_0327_),
    .B(_0267_),
    .C(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2130_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_0318_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2131_ (.I(_0330_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2132_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_0314_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2133_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_1317_),
    .A3(net39),
    .B(_0314_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2134_ (.A1(_0313_),
    .A2(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2135_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_0327_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2136_ (.A1(_0331_),
    .A2(_0333_),
    .B(_0267_),
    .C(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2137_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_0318_),
    .B(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2138_ (.I(_0336_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2139_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2140_ (.I(_0320_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2141_ (.I(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2142_ (.A1(_0317_),
    .A2(_0259_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2143_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_0317_),
    .B(_0313_),
    .C(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2144_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_0333_),
    .B(_0338_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2145_ (.A1(_0337_),
    .A2(_0339_),
    .B1(_0341_),
    .B2(_0342_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2146_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_0259_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2147_ (.A1(_0317_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2148_ (.A1(_0266_),
    .A2(_0312_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2149_ (.I(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2150_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0317_),
    .B1(_0260_),
    .B2(_0344_),
    .C(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2151_ (.I(_0322_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2152_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_0339_),
    .B1(_0348_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2153_ (.A1(_0347_),
    .A2(_0349_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2154_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_0339_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2155_ (.I(_0322_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2156_ (.I(_0345_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2157_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_0351_),
    .B1(_0352_),
    .B2(_0264_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2158_ (.A1(_0350_),
    .A2(_0353_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2159_ (.I(_0346_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2160_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .A2(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2161_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_0339_),
    .B1(_0348_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2162_ (.A1(_0355_),
    .A2(_0356_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2163_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_0321_),
    .B1(_0323_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .C1(_0352_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2164_ (.I(_0357_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2165_ (.I(_0346_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2166_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2167_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_0339_),
    .B1(_0348_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2168_ (.A1(_0359_),
    .A2(_0360_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2169_ (.I(_0345_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2170_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_0321_),
    .B1(_0323_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .C1(_0361_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2171_ (.I(_0362_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2172_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_0358_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2173_ (.I(_0338_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2174_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_0364_),
    .B1(_0348_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2175_ (.A1(_0363_),
    .A2(_0365_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2176_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_0358_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2177_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_0364_),
    .B1(_0348_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2178_ (.A1(_0366_),
    .A2(_0367_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2179_ (.I(_0320_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2180_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_0368_),
    .B1(_0323_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .C1(_0361_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2181_ (.I(_0369_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2182_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_0358_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2183_ (.I(_0322_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2184_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_0364_),
    .B1(_0371_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(_0370_),
    .A2(_0372_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2186_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .A2(_0358_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2187_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_0364_),
    .B1(_0371_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2188_ (.A1(_0373_),
    .A2(_0374_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2189_ (.I(_0345_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2190_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2191_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_0364_),
    .B1(_0371_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2192_ (.A1(_0376_),
    .A2(_0377_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2193_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_0368_),
    .B1(_0323_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .C1(_0361_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2194_ (.I(_0378_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2195_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(_0375_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2196_ (.I(_0338_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2197_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_0380_),
    .B1(_0371_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2198_ (.A1(_0379_),
    .A2(_0381_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2199_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_0375_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2200_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_0380_),
    .B1(_0371_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2201_ (.A1(_0382_),
    .A2(_0383_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2202_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_0375_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2203_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_0380_),
    .B1(_0351_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2204_ (.A1(_0384_),
    .A2(_0385_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2205_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_0375_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2206_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_0380_),
    .B1(_0351_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2207_ (.A1(_0386_),
    .A2(_0387_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2208_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .A2(_0352_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2209_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_0380_),
    .B1(_0351_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2210_ (.A1(_0388_),
    .A2(_0389_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2211_ (.I(_0322_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2212_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_0368_),
    .B1(_0390_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .C1(_0361_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2213_ (.I(_0391_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2214_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0352_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2215_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_0321_),
    .B1(_0351_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2216_ (.A1(_0392_),
    .A2(_0393_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2217_ (.I(_0390_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2218_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0394_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2219_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_0321_),
    .B1(_0352_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2220_ (.A1(_0395_),
    .A2(_0396_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2221_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_0368_),
    .B1(_0390_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .C1(_0361_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2222_ (.I(_0397_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2223_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2224_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2225_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_0318_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2226_ (.A1(_0398_),
    .A2(_0394_),
    .B1(_0354_),
    .B2(_0399_),
    .C(_0400_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2227_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_0368_),
    .B1(_0390_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .C1(_0346_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2228_ (.I(_0401_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2229_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_0338_),
    .B1(_0390_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .C1(_0346_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2230_ (.I(_0402_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2231_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2232_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2233_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_0318_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2234_ (.A1(_0403_),
    .A2(_0394_),
    .B1(_0354_),
    .B2(_0404_),
    .C(_0405_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2235_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2236_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_0267_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2237_ (.A1(_0404_),
    .A2(_0394_),
    .B1(_0354_),
    .B2(_0406_),
    .C(_0407_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2238_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_0267_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2239_ (.A1(_0406_),
    .A2(_0394_),
    .B1(_0354_),
    .B2(_1302_),
    .C(_0408_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2240_ (.A1(_0251_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2241_ (.A1(net12),
    .A2(_1073_),
    .A3(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2242_ (.I(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2243_ (.I(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2244_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2245_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0248_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2246_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0248_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2247_ (.I(_0248_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2248_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2249_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0416_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2250_ (.A1(_0414_),
    .A2(_0415_),
    .A3(_0417_),
    .A4(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2251_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_1079_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2252_ (.I(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2253_ (.A1(_0419_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2254_ (.I(_0416_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2255_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2256_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2257_ (.A1(_0422_),
    .A2(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2258_ (.I(_0416_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2259_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2260_ (.I(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2261_ (.I(_0249_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2262_ (.A1(_0423_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2263_ (.A1(_0430_),
    .A2(\u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2264_ (.I(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2265_ (.A1(_0429_),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2266_ (.A1(_0423_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2267_ (.A1(_0430_),
    .A2(\u_arbiter.i_wb_cpu_rdt[6] ),
    .B(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2268_ (.A1(_0423_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2269_ (.A1(_0430_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2270_ (.A1(_0423_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2271_ (.A1(_1079_),
    .A2(_0337_),
    .B(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2272_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0427_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2273_ (.I0(\u_arbiter.i_wb_cpu_rdt[2] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0427_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2274_ (.A1(_0440_),
    .A2(_0441_),
    .A3(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2275_ (.A1(_0436_),
    .A2(_0438_),
    .A3(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2276_ (.A1(_0248_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2277_ (.A1(_0249_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2278_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2279_ (.A1(_0446_),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2280_ (.A1(_0444_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2281_ (.A1(_0434_),
    .A2(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2282_ (.A1(_0426_),
    .A2(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2283_ (.A1(_0427_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2284_ (.A1(_0430_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2285_ (.I0(\u_arbiter.i_wb_cpu_rdt[1] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_1079_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2286_ (.A1(_0453_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2287_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2288_ (.I(_0447_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2289_ (.A1(_0446_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2290_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_1078_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2291_ (.A1(_0458_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2292_ (.A1(_1078_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2293_ (.A1(_0250_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2294_ (.A1(_0419_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2295_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2296_ (.A1(_0460_),
    .A2(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2297_ (.I(_0446_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2298_ (.I(_0459_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2299_ (.A1(_0466_),
    .A2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(_0465_),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2301_ (.I(_0453_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(_0470_),
    .A2(_0432_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2303_ (.A1(_0429_),
    .A2(_0454_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2304_ (.A1(_0448_),
    .A2(_0471_),
    .B(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2305_ (.I(_0473_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2306_ (.I(_0442_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2307_ (.I(_0410_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2308_ (.I(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2309_ (.A1(_0456_),
    .A2(_0469_),
    .B1(_0474_),
    .B2(_0475_),
    .C(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2310_ (.A1(_0224_),
    .A2(_0413_),
    .B1(_0451_),
    .B2(_0478_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2311_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0416_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2312_ (.I(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2313_ (.A1(_1078_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2314_ (.A1(_0250_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2315_ (.A1(_0480_),
    .A2(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2316_ (.I(_0483_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2317_ (.I(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2318_ (.I(_0440_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2319_ (.I(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2320_ (.A1(_0456_),
    .A2(_0485_),
    .B1(_0474_),
    .B2(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2321_ (.I(_0411_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2322_ (.A1(_0222_),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2323_ (.A1(_0413_),
    .A2(_0488_),
    .B(_0490_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2324_ (.I(_0470_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2325_ (.A1(_1078_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2326_ (.A1(_0250_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2327_ (.A1(_0446_),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2328_ (.A1(_0484_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2329_ (.I(_0473_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2330_ (.A1(_0476_),
    .A2(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2331_ (.I(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2332_ (.A1(_0491_),
    .A2(_0495_),
    .B(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2333_ (.I(_0493_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2334_ (.A1(_0500_),
    .A2(_0444_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2335_ (.I(_0480_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2336_ (.A1(_0470_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2337_ (.A1(_0426_),
    .A2(_0433_),
    .A3(_0501_),
    .B(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2338_ (.I(_0411_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2339_ (.A1(_0480_),
    .A2(_0493_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2340_ (.A1(_0428_),
    .A2(_0454_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2341_ (.A1(_0453_),
    .A2(_0432_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2342_ (.A1(_0506_),
    .A2(_0507_),
    .B(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2343_ (.A1(_0410_),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2344_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2345_ (.A1(_1320_),
    .A2(_0505_),
    .B1(_0441_),
    .B2(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2346_ (.A1(_0499_),
    .A2(_0504_),
    .B(_0512_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2347_ (.I(_0253_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2348_ (.I(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2349_ (.I(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2350_ (.A1(_0429_),
    .A2(_0432_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2351_ (.I(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2352_ (.A1(_0448_),
    .A2(_0459_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2353_ (.I(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2354_ (.A1(_1079_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2355_ (.A1(_0430_),
    .A2(\u_arbiter.i_wb_cpu_rdt[11] ),
    .B(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2356_ (.A1(_0427_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2357_ (.A1(_0250_),
    .A2(\u_arbiter.i_wb_cpu_rdt[10] ),
    .B(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2358_ (.I(_0523_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2359_ (.A1(_0521_),
    .A2(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2360_ (.A1(_0519_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2361_ (.A1(_0465_),
    .A2(_0495_),
    .A3(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2362_ (.I(_0500_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2363_ (.I(_0473_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2364_ (.I(_0411_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2365_ (.A1(_0491_),
    .A2(_0528_),
    .B1(_0438_),
    .B2(_0529_),
    .C(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2366_ (.A1(_0517_),
    .A2(_0527_),
    .B(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2367_ (.A1(_1209_),
    .A2(_0515_),
    .B(_0532_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2368_ (.I(_0429_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2369_ (.A1(_0502_),
    .A2(_0457_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2370_ (.A1(_0468_),
    .A2(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2371_ (.A1(_0513_),
    .A2(_0509_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2372_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2373_ (.A1(_0533_),
    .A2(_0535_),
    .B(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2374_ (.I(_0436_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2375_ (.A1(_1266_),
    .A2(_0514_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2376_ (.A1(_0450_),
    .A2(_0538_),
    .B1(_0511_),
    .B2(_0539_),
    .C(_0540_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2377_ (.I(_1235_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2378_ (.I(_0513_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2379_ (.A1(_0460_),
    .A2(_0463_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2380_ (.I(_0494_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2381_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_1080_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2382_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_1080_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2383_ (.A1(_0545_),
    .A2(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2384_ (.I(_0506_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2385_ (.A1(_0548_),
    .A2(_0482_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2386_ (.A1(_0525_),
    .A2(_0547_),
    .B(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2387_ (.A1(_0475_),
    .A2(_0543_),
    .B1(_0544_),
    .B2(_0467_),
    .C(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2388_ (.I(_0424_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2389_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2390_ (.I(_0516_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2391_ (.A1(_0554_),
    .A2(_0468_),
    .B(_0509_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2392_ (.A1(_0479_),
    .A2(_0457_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2393_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2394_ (.A1(_0553_),
    .A2(_0555_),
    .B1(_0557_),
    .B2(_0434_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2395_ (.A1(_0517_),
    .A2(_0551_),
    .B(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2396_ (.A1(_0542_),
    .A2(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2397_ (.A1(_0541_),
    .A2(_0515_),
    .B(_0560_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2398_ (.I(_0509_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2399_ (.I(_0521_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2400_ (.A1(_0415_),
    .A2(_0539_),
    .B(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2401_ (.A1(_0552_),
    .A2(_0483_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2402_ (.A1(_0486_),
    .A2(_0543_),
    .B1(_0519_),
    .B2(_0563_),
    .C(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2403_ (.A1(_0517_),
    .A2(_0565_),
    .B(_0503_),
    .C(_0561_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2404_ (.A1(_0467_),
    .A2(_0561_),
    .B(_0566_),
    .C(_0514_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2405_ (.A1(_0215_),
    .A2(_0515_),
    .B(_0567_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2406_ (.I(_0254_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2407_ (.A1(_0539_),
    .A2(_0438_),
    .A3(_0525_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2408_ (.A1(_0441_),
    .A2(_0543_),
    .B1(_0519_),
    .B2(_0569_),
    .C(_0564_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2409_ (.A1(_0466_),
    .A2(_0472_),
    .B1(_0570_),
    .B2(_0517_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2410_ (.A1(_0568_),
    .A2(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2411_ (.A1(_1029_),
    .A2(_0515_),
    .B(_0572_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2412_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_1082_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2413_ (.A1(_0475_),
    .A2(_0482_),
    .A3(_0534_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2414_ (.A1(_0424_),
    .A2(_0543_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2415_ (.A1(_0564_),
    .A2(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2416_ (.A1(_0533_),
    .A2(_0574_),
    .A3(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2417_ (.I(_0480_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2418_ (.I(_0493_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2419_ (.A1(_0578_),
    .A2(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2420_ (.A1(_0426_),
    .A2(_0449_),
    .B1(_0580_),
    .B2(_0442_),
    .C(_0433_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2421_ (.I(_0494_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2422_ (.I(_0471_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2423_ (.A1(_0442_),
    .A2(_0582_),
    .B(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2424_ (.A1(_0530_),
    .A2(_0508_),
    .A3(_0581_),
    .A4(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2425_ (.A1(_0510_),
    .A2(_0573_),
    .B1(_0577_),
    .B2(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2426_ (.A1(_1039_),
    .A2(_0515_),
    .B(_0586_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2427_ (.I(_0514_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2428_ (.I(_0510_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2429_ (.I(_1081_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2430_ (.I(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2431_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2432_ (.I(_0454_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2433_ (.A1(_0500_),
    .A2(_0482_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2434_ (.A1(_0502_),
    .A2(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2435_ (.A1(_0486_),
    .A2(_0594_),
    .B(_0575_),
    .C(_0470_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2436_ (.A1(_0491_),
    .A2(_0486_),
    .A3(_0580_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2437_ (.A1(_0592_),
    .A2(_0595_),
    .B(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2438_ (.I(_0507_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2439_ (.A1(_0487_),
    .A2(_0544_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2440_ (.A1(_0598_),
    .A2(_0599_),
    .B(_0536_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2441_ (.A1(_0588_),
    .A2(_0591_),
    .B1(_0597_),
    .B2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2442_ (.A1(_1040_),
    .A2(_0587_),
    .B(_0601_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2443_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_1081_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(_0471_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2445_ (.A1(_1080_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2446_ (.A1(_0251_),
    .A2(\u_arbiter.i_wb_cpu_rdt[4] ),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2447_ (.A1(_0455_),
    .A2(_0575_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2448_ (.A1(_0575_),
    .A2(_0594_),
    .B(_0455_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2449_ (.A1(_0453_),
    .A2(_0454_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2450_ (.A1(_0605_),
    .A2(_0606_),
    .B1(_0607_),
    .B2(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2451_ (.I(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2452_ (.A1(_0441_),
    .A2(_0582_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2453_ (.A1(_0579_),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0602_),
    .C(_0583_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2454_ (.A1(_0603_),
    .A2(_0610_),
    .B1(_0611_),
    .B2(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2455_ (.A1(_0588_),
    .A2(_0602_),
    .B1(_0613_),
    .B2(_0498_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2456_ (.A1(_1245_),
    .A2(_0587_),
    .B(_0614_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2457_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_0413_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2458_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_0589_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2459_ (.A1(_0482_),
    .A2(_0556_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2460_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2461_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2462_ (.A1(_0553_),
    .A2(_0619_),
    .B(_0456_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2463_ (.I(_0418_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2465_ (.A1(_0552_),
    .A2(_0502_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2466_ (.A1(_0414_),
    .A2(_0523_),
    .A3(_0424_),
    .A4(_0518_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2467_ (.I(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2468_ (.A1(_0593_),
    .A2(_0623_),
    .B(_0625_),
    .C(_0618_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2469_ (.A1(_0552_),
    .A2(_0463_),
    .B(_0459_),
    .C(_0458_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2470_ (.A1(_0438_),
    .A2(_0464_),
    .B(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2471_ (.A1(_0626_),
    .A2(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2472_ (.A1(_0622_),
    .A2(_0485_),
    .B1(_0544_),
    .B2(_0546_),
    .C(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_0458_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2474_ (.A1(_0475_),
    .A2(_0631_),
    .B1(_0582_),
    .B2(_0621_),
    .C(_0433_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2475_ (.A1(_0620_),
    .A2(_0630_),
    .B1(_0632_),
    .B2(_0533_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2476_ (.A1(_0466_),
    .A2(_0500_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _2477_ (.A1(_0466_),
    .A2(_0546_),
    .B1(_0448_),
    .B2(_0616_),
    .C1(_0634_),
    .C2(_0622_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2478_ (.A1(_0598_),
    .A2(_0635_),
    .B(_0537_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2479_ (.A1(_0588_),
    .A2(_0616_),
    .B1(_0633_),
    .B2(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(_0615_),
    .A2(_0637_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2481_ (.I(_0411_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2482_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2483_ (.A1(_0297_),
    .A2(_1209_),
    .A3(_1034_),
    .B(_1232_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2484_ (.A1(_0476_),
    .A2(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2485_ (.I(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2487_ (.A1(_0639_),
    .A2(_0642_),
    .B(_0643_),
    .C(_0586_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2488_ (.I(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2489_ (.A1(_0644_),
    .A2(_0640_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2490_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_0640_),
    .B(_0645_),
    .C(_0489_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2491_ (.A1(_0601_),
    .A2(_0646_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2492_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2493_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0640_),
    .B(_0638_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2494_ (.A1(_0647_),
    .A2(_0642_),
    .B1(_0648_),
    .B2(_0614_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2495_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_1081_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2496_ (.A1(_0608_),
    .A2(_0607_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2497_ (.A1(_0425_),
    .A2(_0543_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2498_ (.A1(_0526_),
    .A2(_0651_),
    .B(_0607_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2499_ (.A1(_0546_),
    .A2(_0650_),
    .B(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(_0524_),
    .A2(_0579_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2501_ (.A1(_0578_),
    .A2(_0649_),
    .B(_0654_),
    .C(_0634_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2502_ (.I(_0471_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2503_ (.A1(_0546_),
    .A2(_0557_),
    .B(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2504_ (.A1(_0583_),
    .A2(_0653_),
    .B1(_0655_),
    .B2(_0657_),
    .C(_0496_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2505_ (.A1(_0474_),
    .A2(_0649_),
    .B(_0658_),
    .C(_0477_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2506_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_0568_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0642_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2508_ (.A1(_0642_),
    .A2(_0659_),
    .A3(_0660_),
    .B(_0661_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2509_ (.A1(_0414_),
    .A2(_0485_),
    .B(_0491_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2510_ (.A1(_0539_),
    .A2(_0527_),
    .B(_0651_),
    .C(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2511_ (.I(_0506_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2512_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_1082_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2513_ (.A1(_0414_),
    .A2(_0528_),
    .B1(_0664_),
    .B2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2514_ (.A1(_0592_),
    .A2(_0539_),
    .B1(_0598_),
    .B2(_0666_),
    .C(_0508_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2515_ (.A1(_0498_),
    .A2(_0663_),
    .A3(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2516_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0476_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2517_ (.A1(_0641_),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2518_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_0641_),
    .B1(_0665_),
    .B2(_0588_),
    .C(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2519_ (.A1(_0668_),
    .A2(_0671_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2520_ (.A1(_0467_),
    .A2(_0464_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2521_ (.A1(_0495_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2522_ (.A1(_0475_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2523_ (.I(_0593_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2524_ (.A1(_0553_),
    .A2(_0675_),
    .B(_0624_),
    .C(_0575_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2525_ (.A1(_0533_),
    .A2(_0674_),
    .A3(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2526_ (.A1(_0553_),
    .A2(_0533_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2527_ (.A1(_0592_),
    .A2(_0503_),
    .B(_0678_),
    .C(_0529_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2528_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .S(_0590_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2529_ (.A1(_0677_),
    .A2(_0679_),
    .B1(_0680_),
    .B2(_0474_),
    .C(_0477_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2530_ (.A1(_1320_),
    .A2(_1265_),
    .A3(_1204_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2531_ (.A1(_0297_),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2532_ (.A1(_1232_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2533_ (.A1(_0530_),
    .A2(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2534_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_0542_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2535_ (.A1(_0297_),
    .A2(_0682_),
    .B(_0218_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2536_ (.A1(_0254_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2537_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2538_ (.A1(_0681_),
    .A2(_0686_),
    .B(_0689_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2539_ (.A1(_0254_),
    .A2(_0684_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2540_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_0688_),
    .B1(_0690_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(_0637_),
    .A2(_0691_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2542_ (.A1(_0487_),
    .A2(_0631_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2543_ (.A1(_0545_),
    .A2(_0535_),
    .B(_0491_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2544_ (.A1(_0672_),
    .A2(_0692_),
    .B(_0693_),
    .C(_0676_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2545_ (.I(_0420_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2546_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_1082_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2547_ (.A1(_0695_),
    .A2(_0557_),
    .B1(_0696_),
    .B2(_0664_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2548_ (.A1(_0420_),
    .A2(_0494_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2549_ (.A1(_0487_),
    .A2(_0631_),
    .B(_0433_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2550_ (.A1(_0598_),
    .A2(_0697_),
    .B1(_0698_),
    .B2(_0699_),
    .C(_0537_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2551_ (.A1(_0694_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2552_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_0688_),
    .B1(_0690_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_0696_),
    .C2(_0588_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2553_ (.A1(_0701_),
    .A2(_0702_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2554_ (.I(_0417_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2555_ (.A1(_0605_),
    .A2(_0464_),
    .B(_0627_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2556_ (.A1(_0626_),
    .A2(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2557_ (.A1(_0703_),
    .A2(_0484_),
    .B1(_0544_),
    .B2(_0553_),
    .C(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2558_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .S(_0589_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2559_ (.A1(_0703_),
    .A2(_0557_),
    .B1(_0707_),
    .B2(_0664_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2560_ (.A1(_0620_),
    .A2(_0706_),
    .B1(_0708_),
    .B2(_0603_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2561_ (.A1(_0537_),
    .A2(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2562_ (.A1(_0476_),
    .A2(_0687_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2563_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_0685_),
    .B1(_0711_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2564_ (.A1(_0477_),
    .A2(_0561_),
    .A3(_0707_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2565_ (.A1(_0710_),
    .A2(_0712_),
    .A3(_0713_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2566_ (.A1(_0589_),
    .A2(\u_arbiter.i_wb_cpu_rdt[29] ),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2567_ (.A1(_0251_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2568_ (.A1(_0457_),
    .A2(_0715_),
    .B(_0583_),
    .C(_0578_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2569_ (.A1(_0415_),
    .A2(_0485_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2570_ (.A1(_0618_),
    .A2(_0623_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2571_ (.A1(_0624_),
    .A2(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2572_ (.A1(_0717_),
    .A2(_0719_),
    .B(_0620_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2573_ (.A1(_0654_),
    .A2(_0716_),
    .B(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2574_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_0685_),
    .B1(_0711_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2575_ (.A1(_0511_),
    .A2(_0715_),
    .B1(_0721_),
    .B2(_0498_),
    .C(_0722_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2576_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_0590_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2577_ (.A1(_0524_),
    .A2(_0425_),
    .B(_0562_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2578_ (.A1(_0562_),
    .A2(_0524_),
    .B1(_0569_),
    .B2(_0724_),
    .C(_0549_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2579_ (.A1(_0695_),
    .A2(_0485_),
    .B(_0718_),
    .C(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2580_ (.A1(_0620_),
    .A2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2581_ (.A1(_0510_),
    .A2(_0723_),
    .B1(_0727_),
    .B2(_0514_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2582_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_0688_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2583_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2584_ (.A1(_1320_),
    .A2(_0297_),
    .B(_0222_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2585_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_1222_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2586_ (.A1(_0732_),
    .A2(_0731_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2587_ (.A1(_0730_),
    .A2(_0731_),
    .B(_0733_),
    .C(_0225_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2588_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_0225_),
    .B(_0690_),
    .C(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2589_ (.A1(_0728_),
    .A2(_0729_),
    .A3(_0735_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2590_ (.A1(_0419_),
    .A2(_0421_),
    .B(_0425_),
    .C(_0449_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2591_ (.A1(_0621_),
    .A2(_0501_),
    .A3(_0534_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2592_ (.A1(_0592_),
    .A2(_0736_),
    .A3(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2593_ (.A1(_1080_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2594_ (.A1(_0251_),
    .A2(\u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2595_ (.A1(_0459_),
    .A2(_0634_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2596_ (.A1(_0425_),
    .A2(_0582_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2597_ (.A1(_0740_),
    .A2(_0502_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2598_ (.A1(_0621_),
    .A2(_0519_),
    .B1(_0743_),
    .B2(_0579_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2599_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0742_),
    .B2(_0744_),
    .C(_0554_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2600_ (.A1(_0470_),
    .A2(_0738_),
    .B(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2601_ (.A1(_0579_),
    .A2(_0442_),
    .B1(_0548_),
    .B2(_0621_),
    .C(_0583_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2602_ (.A1(_0746_),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2603_ (.A1(_0622_),
    .A2(_0510_),
    .B1(_0748_),
    .B2(_0497_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2604_ (.A1(_0218_),
    .A2(_0732_),
    .B(_0638_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2605_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_0542_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2606_ (.A1(_0749_),
    .A2(_0750_),
    .B1(_0751_),
    .B2(_0219_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2607_ (.A1(_1310_),
    .A2(_0222_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2608_ (.A1(_1222_),
    .A2(_1292_),
    .A3(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2609_ (.A1(_1232_),
    .A2(_0753_),
    .B(_0513_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2610_ (.I(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2611_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2612_ (.I(_0754_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2613_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_0505_),
    .B(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2614_ (.A1(_0730_),
    .A2(_0756_),
    .B1(_0758_),
    .B2(_0586_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2615_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2616_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_0505_),
    .B(_0757_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2617_ (.A1(_0759_),
    .A2(_0756_),
    .B1(_0760_),
    .B2(_0560_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2618_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2619_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_0505_),
    .B(_0757_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2620_ (.A1(_0761_),
    .A2(_0756_),
    .B1(_0762_),
    .B2(_0567_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2621_ (.I(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2622_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_0505_),
    .B(_0757_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2623_ (.A1(_0763_),
    .A2(_0756_),
    .B1(_0764_),
    .B2(_0572_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2624_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2625_ (.A1(_0552_),
    .A2(_0483_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2626_ (.A1(_0438_),
    .A2(_0465_),
    .B(_0766_),
    .C(_0619_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2627_ (.A1(_0622_),
    .A2(_0619_),
    .B(_0767_),
    .C(_0456_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2628_ (.A1(_0656_),
    .A2(_0557_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2629_ (.A1(_0417_),
    .A2(_0617_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2630_ (.A1(_0516_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2631_ (.A1(_0500_),
    .A2(_0483_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2632_ (.A1(_0424_),
    .A2(_0493_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2633_ (.A1(_0444_),
    .A2(_0773_),
    .B(_0608_),
    .C(_0480_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2634_ (.A1(_0771_),
    .A2(_0772_),
    .B(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2635_ (.I(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2636_ (.A1(_0769_),
    .A2(_0743_),
    .B1(_0776_),
    .B2(_0622_),
    .C(_0496_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2637_ (.A1(_0528_),
    .A2(_0508_),
    .B1(_0768_),
    .B2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2638_ (.A1(_0542_),
    .A2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2639_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0489_),
    .B(_0755_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2640_ (.A1(_0765_),
    .A2(_0756_),
    .B1(_0779_),
    .B2(_0780_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2641_ (.I(_0757_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2642_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_0589_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2643_ (.A1(_0548_),
    .A2(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2644_ (.A1(_0421_),
    .A2(_0578_),
    .B(_0656_),
    .C(_0556_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2645_ (.A1(_0545_),
    .A2(_0464_),
    .B(_0467_),
    .C(_0458_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2646_ (.A1(_0420_),
    .A2(_0519_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2647_ (.A1(_0766_),
    .A2(_0618_),
    .A3(_0698_),
    .A4(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2648_ (.A1(_0462_),
    .A2(_0741_),
    .B1(_0785_),
    .B2(_0787_),
    .C(_0554_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2649_ (.A1(_0444_),
    .A2(_0773_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2650_ (.A1(_0421_),
    .A2(_0434_),
    .A3(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2651_ (.A1(_0656_),
    .A2(_0503_),
    .A3(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2652_ (.A1(_0788_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2653_ (.A1(_0783_),
    .A2(_0784_),
    .B(_0496_),
    .C(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2654_ (.A1(_0474_),
    .A2(_0782_),
    .B(_0793_),
    .C(_0477_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2655_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0568_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2656_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0781_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2657_ (.A1(_0781_),
    .A2(_0794_),
    .A3(_0795_),
    .B(_0796_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2658_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .S(_1081_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(_0576_),
    .A2(_0618_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2660_ (.I(_0507_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2661_ (.A1(_0417_),
    .A2(_0776_),
    .B1(_0798_),
    .B2(_0771_),
    .C(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2662_ (.A1(_0703_),
    .A2(_0578_),
    .B1(_0548_),
    .B2(_0797_),
    .C(_0656_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2663_ (.A1(_0529_),
    .A2(_0800_),
    .A3(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2664_ (.A1(_0529_),
    .A2(_0797_),
    .B(_0802_),
    .C(_0412_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2665_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0568_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2666_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0755_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2667_ (.A1(_0781_),
    .A2(_0803_),
    .A3(_0804_),
    .B(_0805_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2668_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .S(_0590_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2669_ (.A1(_0631_),
    .A2(_0484_),
    .B(_0576_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2670_ (.A1(_0524_),
    .A2(_0741_),
    .B(_0554_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2671_ (.A1(_0415_),
    .A2(_0774_),
    .B1(_0807_),
    .B2(_0808_),
    .C(_0799_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2672_ (.A1(_0466_),
    .A2(_0799_),
    .B(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2673_ (.A1(_0529_),
    .A2(_0806_),
    .B(_0810_),
    .C(_0412_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2674_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0568_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2675_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0755_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2676_ (.A1(_0781_),
    .A2(_0811_),
    .A3(_0812_),
    .B(_0813_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2677_ (.A1(_0562_),
    .A2(_0619_),
    .B(_0576_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2678_ (.A1(_1082_),
    .A2(_0337_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2679_ (.A1(_0590_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_0496_),
    .C(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2680_ (.A1(_0254_),
    .A2(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2681_ (.A1(_0414_),
    .A2(_0774_),
    .B1(_0814_),
    .B2(_0456_),
    .C(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2682_ (.A1(_1033_),
    .A2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2683_ (.A1(_0530_),
    .A2(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2684_ (.A1(_1266_),
    .A2(_0732_),
    .B(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0755_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2686_ (.A1(_0781_),
    .A2(_0818_),
    .A3(_0821_),
    .B(_0822_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2687_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_1083_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2688_ (.A1(_0766_),
    .A2(_0719_),
    .B(_0620_),
    .C(_0530_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2689_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_0489_),
    .B1(_0511_),
    .B2(_0823_),
    .C(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2690_ (.I(_0825_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2691_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2692_ (.A1(_0277_),
    .A2(_0243_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2693_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2694_ (.A1(_0826_),
    .A2(_0827_),
    .B(_0828_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2695_ (.I0(\u_cpu.cpu.alu.cmp_r ),
    .I1(_0304_),
    .S(_1232_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2696_ (.I(_0829_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2697_ (.I(_1288_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2698_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2699_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_0832_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2701_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_0831_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2702_ (.I(_0833_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2703_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_0831_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2704_ (.I(_0834_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2705_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_0831_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2706_ (.I(_0835_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2707_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_0831_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2708_ (.I(_0836_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2709_ (.I(_0830_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2710_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2711_ (.I(_0838_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2712_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_0837_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2713_ (.I(_0839_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2714_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_0837_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2715_ (.I(_0840_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2716_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_0837_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2717_ (.I(_0841_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2718_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_0837_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2719_ (.I(_0842_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2720_ (.I(_1288_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2721_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2722_ (.I(_0844_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2723_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_0843_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2724_ (.I(_0845_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2725_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_0843_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2726_ (.I(_0846_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2727_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_0843_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2728_ (.I(_0847_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2729_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_0843_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2730_ (.I(_0848_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2731_ (.I(_1288_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2732_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2733_ (.I(_0850_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2734_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_0849_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2735_ (.I(_0851_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2736_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_0849_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2737_ (.I(_0852_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2738_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_0849_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2739_ (.I(_0853_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2740_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_0849_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2741_ (.I(_0854_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2742_ (.I(_1288_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2743_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2744_ (.I(_0856_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2745_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_0855_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2746_ (.I(_0857_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2747_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_0855_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2748_ (.I(_0858_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2749_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_0855_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2750_ (.I(_0859_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2751_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_0855_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2752_ (.I(_0860_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2753_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_0830_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2754_ (.I(_0861_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2755_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_0830_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2756_ (.I(_0862_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2757_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_0830_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2758_ (.I(_0863_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2759_ (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2760_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_0233_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2761_ (.A1(_0864_),
    .A2(_0233_),
    .B(_0865_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2762_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_0243_),
    .B(_0233_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2763_ (.A1(_0228_),
    .A2(_0231_),
    .B(_0243_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2764_ (.A1(_0228_),
    .A2(_0231_),
    .B(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2765_ (.A1(_0864_),
    .A2(_0866_),
    .B1(_0868_),
    .B2(_0233_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2766_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(_1281_),
    .B(_1247_),
    .C(_0257_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2767_ (.A1(_1279_),
    .A2(_0257_),
    .B(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2768_ (.A1(_1026_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2769_ (.A1(_1267_),
    .A2(_0870_),
    .B(_0871_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2770_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_0243_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2771_ (.A1(_0868_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2772_ (.A1(_0870_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2773_ (.A1(_0216_),
    .A2(_0870_),
    .B(_0874_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2774_ (.A1(_1231_),
    .A2(_0237_),
    .B(net2),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2775_ (.I(_0875_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2776_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2777_ (.A1(net2),
    .A2(_0238_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2778_ (.I(_0878_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2779_ (.I(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2780_ (.A1(_1071_),
    .A2(_0877_),
    .B1(_0880_),
    .B2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2781_ (.I(_0881_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2782_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0877_),
    .B1(_0880_),
    .B2(_1084_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2783_ (.I(_0882_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2784_ (.A1(_1084_),
    .A2(_0877_),
    .B1(_0880_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2785_ (.I(_0883_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2786_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0877_),
    .B1(_0880_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2787_ (.I(_0884_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2788_ (.I(_0876_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2789_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0885_),
    .B1(_0880_),
    .B2(_1100_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2790_ (.I(_0886_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2791_ (.I(_0879_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2792_ (.A1(_1100_),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2793_ (.I(_0888_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2794_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2795_ (.I(_0889_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2796_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2797_ (.I(_0890_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2798_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2799_ (.I(_0891_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2800_ (.I(_0875_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2801_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0892_),
    .B1(_0887_),
    .B2(_1124_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2802_ (.I(_0893_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2803_ (.I(_0879_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2804_ (.A1(_1124_),
    .A2(_0892_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2805_ (.I(_0895_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2806_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_0892_),
    .B1(_0894_),
    .B2(_1133_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2807_ (.I(_0896_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2808_ (.A1(_1133_),
    .A2(_0892_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2809_ (.I(_0897_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2810_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_0892_),
    .B1(_0894_),
    .B2(_1140_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2811_ (.I(_0898_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2812_ (.I(_0875_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2813_ (.A1(_1140_),
    .A2(_0899_),
    .B1(_0894_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2814_ (.I(_0900_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2815_ (.I(_0879_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2816_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(_1147_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2817_ (.I(_0902_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2818_ (.A1(_1147_),
    .A2(_0899_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2819_ (.I(_0903_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2820_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2821_ (.I(_0904_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2822_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0899_),
    .B1(_0901_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2823_ (.I(_0905_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2824_ (.I(_0875_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2825_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_0906_),
    .B1(_0901_),
    .B2(_1160_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(_0907_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2827_ (.I(_0878_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2828_ (.A1(_1160_),
    .A2(_0906_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2829_ (.I(_0909_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2830_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0906_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2831_ (.I(_0910_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2832_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0906_),
    .B1(_0908_),
    .B2(_1169_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2833_ (.I(_0911_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2834_ (.A1(_1169_),
    .A2(_0906_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2835_ (.I(_0912_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2836_ (.I(_0875_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2837_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_0913_),
    .B1(_0908_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2838_ (.I(_0914_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2839_ (.I(_0878_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2840_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0913_),
    .B1(_0915_),
    .B2(_1181_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2841_ (.I(_0916_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2842_ (.A1(_1181_),
    .A2(_0913_),
    .B1(_0915_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2843_ (.I(_0917_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2844_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_0913_),
    .B1(_0915_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2845_ (.I(_0918_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2846_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0913_),
    .B1(_0915_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2847_ (.I(_0919_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2848_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0876_),
    .B1(_0915_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2849_ (.I(_0920_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2850_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_0876_),
    .B1(_0879_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2851_ (.I(_0921_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2852_ (.A1(_1040_),
    .A2(_1049_),
    .A3(_1042_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2853_ (.A1(_1052_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2854_ (.I(_1327_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2855_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2856_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_1296_),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2857_ (.A1(_0923_),
    .A2(_1307_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2858_ (.A1(_0923_),
    .A2(_0926_),
    .B1(_0927_),
    .B2(_1243_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2859_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0876_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2860_ (.A1(_0246_),
    .A2(_0238_),
    .A3(_0928_),
    .B(_0929_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2861_ (.A1(_0218_),
    .A2(_0242_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2862_ (.A1(_0513_),
    .A2(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2863_ (.I(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2864_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0638_),
    .B(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2865_ (.A1(_1218_),
    .A2(_0932_),
    .B1(_0933_),
    .B2(_0749_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2866_ (.A1(_0695_),
    .A2(_0434_),
    .A3(_0501_),
    .A4(_0534_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2867_ (.A1(_0421_),
    .A2(_0631_),
    .B1(_0582_),
    .B2(_0486_),
    .C(_0741_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2868_ (.A1(_0462_),
    .A2(_0741_),
    .B1(_0786_),
    .B2(_0935_),
    .C(_0554_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_0799_),
    .A2(_0936_),
    .B(_0561_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2870_ (.A1(_0528_),
    .A2(_0487_),
    .B1(_0664_),
    .B2(_0695_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2871_ (.A1(_0934_),
    .A2(_0937_),
    .B1(_0938_),
    .B2(_0598_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2872_ (.A1(_0587_),
    .A2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2873_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0930_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2874_ (.A1(_1386_),
    .A2(_0930_),
    .B(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2875_ (.A1(_0695_),
    .A2(_0511_),
    .B1(_0942_),
    .B2(_0489_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2876_ (.A1(_0940_),
    .A2(_0943_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2877_ (.A1(_0528_),
    .A2(_0441_),
    .B1(_0544_),
    .B2(_0545_),
    .C1(_0664_),
    .C2(_0703_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2878_ (.A1(_0417_),
    .A2(_0495_),
    .A3(_0634_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2879_ (.A1(_0611_),
    .A2(_0619_),
    .A3(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2880_ (.A1(_0771_),
    .A2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2881_ (.A1(_0603_),
    .A2(_0944_),
    .B(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2882_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0638_),
    .B1(_0498_),
    .B2(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2883_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_0932_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2884_ (.A1(_0608_),
    .A2(_0449_),
    .B(_0509_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2885_ (.A1(_0542_),
    .A2(_0703_),
    .A3(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2886_ (.A1(_0932_),
    .A2(_0949_),
    .B(_0950_),
    .C(_0952_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2887_ (.A1(_1389_),
    .A2(_0930_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2888_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0930_),
    .B(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2889_ (.A1(_0592_),
    .A2(_0484_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2890_ (.A1(_0799_),
    .A2(_0951_),
    .A3(_0955_),
    .B(_0415_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2891_ (.A1(_0457_),
    .A2(_0603_),
    .B1(_0549_),
    .B2(_0517_),
    .C(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2892_ (.A1(_0587_),
    .A2(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2893_ (.A1(_0587_),
    .A2(_0954_),
    .B(_0958_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2894_ (.A1(_0429_),
    .A2(_0580_),
    .A3(_0593_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2895_ (.A1(_0501_),
    .A2(_0603_),
    .A3(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2896_ (.A1(_0561_),
    .A2(_0534_),
    .A3(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2897_ (.A1(_0412_),
    .A2(_0562_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2898_ (.A1(_0961_),
    .A2(_0962_),
    .B(_0931_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2899_ (.A1(_1389_),
    .A2(_0932_),
    .B1(_0963_),
    .B2(_0669_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2900_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_0413_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2901_ (.A1(_0728_),
    .A2(_0964_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2902_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(\u_arbiter.o_wb_cpu_adr[1] ),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2903_ (.A1(_1083_),
    .A2(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2904_ (.A1(_0247_),
    .A2(_0966_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2905_ (.I(_0252_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2906_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2907_ (.I(_0968_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2908_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_0967_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2909_ (.I(_0969_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2910_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0967_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2911_ (.I(_0970_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2912_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_0967_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2913_ (.I(_0971_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2914_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0967_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2915_ (.I(_0972_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2916_ (.I(_0252_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2917_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2918_ (.I(_0974_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2919_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_0973_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2920_ (.I(_0975_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2921_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0973_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2922_ (.I(_0976_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2923_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_0973_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2924_ (.I(_0977_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2925_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0973_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2926_ (.I(_0978_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2927_ (.I(_0252_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2928_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2929_ (.I(_0980_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2930_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0979_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2931_ (.I(_0981_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2932_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0979_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2933_ (.I(_0982_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2934_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_0979_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2935_ (.I(_0983_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2936_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0979_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2937_ (.I(_0984_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2938_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_0252_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2939_ (.I(_0985_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2940_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2941_ (.A1(_1045_),
    .A2(_0986_),
    .B(_1051_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2942_ (.A1(_0277_),
    .A2(_1052_),
    .B1(_1254_),
    .B2(_1247_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2943_ (.I(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2944_ (.I0(_0987_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .S(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2945_ (.I(_0990_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2946_ (.A1(_1033_),
    .A2(_1204_),
    .B1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .B2(_1046_),
    .C(_0988_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2947_ (.A1(_0986_),
    .A2(_0989_),
    .B1(_0991_),
    .B2(_1051_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2948_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2949_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2950_ (.A1(_0993_),
    .A2(_1262_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2951_ (.A1(_1047_),
    .A2(_1033_),
    .A3(_0988_),
    .A4(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2952_ (.A1(_0992_),
    .A2(_0989_),
    .B(_0995_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2953_ (.A1(_1039_),
    .A2(_1050_),
    .B(_0989_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2954_ (.A1(_0993_),
    .A2(_0989_),
    .B1(_0996_),
    .B2(_1261_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2955_ (.I(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2956_ (.A1(_0277_),
    .A2(_1253_),
    .B(_1262_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2957_ (.A1(_1047_),
    .A2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2958_ (.A1(_0997_),
    .A2(_0998_),
    .B1(_0999_),
    .B2(_1261_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2959_ (.A1(_0277_),
    .A2(_1262_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2960_ (.I0(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .I1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .S(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2961_ (.I(_1001_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2962_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2963_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(_1246_),
    .A3(_1315_),
    .A4(_1245_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2964_ (.A1(_1248_),
    .A2(_0281_),
    .A3(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2965_ (.A1(_1260_),
    .A2(_1004_),
    .B(_0282_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2966_ (.A1(_1002_),
    .A2(_1004_),
    .B(_1005_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2967_ (.A1(_0922_),
    .A2(_1260_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2968_ (.A1(_0922_),
    .A2(_1249_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2969_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_1038_),
    .B(_1234_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2970_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_1000_),
    .A3(_1007_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2971_ (.A1(_1006_),
    .A2(_1007_),
    .A3(_1008_),
    .B(_1009_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2972_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_0413_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2973_ (.A1(_0537_),
    .A2(_1010_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2974_ (.A1(_1047_),
    .A2(_0287_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2975_ (.A1(_0246_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_0828_),
    .B(_1011_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2976_ (.A1(_0412_),
    .A2(_0286_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2977_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2978_ (.A1(_0877_),
    .A2(_1012_),
    .B(_1013_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2979_ (.A1(_1353_),
    .A2(_0024_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2980_ (.A1(_1214_),
    .A2(_1014_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2981_ (.A1(_1027_),
    .A2(_1014_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2982_ (.A1(_0282_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2983_ (.I(_1015_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2984_ (.A1(_1020_),
    .A2(_1022_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2985_ (.A1(_0271_),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2986_ (.A1(_1016_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2987_ (.A1(_0255_),
    .A2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2988_ (.A1(_0269_),
    .A2(_1019_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2989_ (.D(_0027_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2990_ (.D(_0028_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2991_ (.D(_0029_),
    .CLK(net65),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2992_ (.D(_0030_),
    .CLK(net65),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2993_ (.D(_0031_),
    .CLK(net66),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2994_ (.D(_0007_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2995_ (.D(_0008_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2996_ (.D(_0009_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2997_ (.D(_0010_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2998_ (.D(_0011_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2999_ (.D(_0012_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3000_ (.D(_0000_),
    .CLK(net65),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3001_ (.D(_0001_),
    .CLK(net65),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3002_ (.D(_0002_),
    .CLK(net65),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3003_ (.D(_0003_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3004_ (.D(_0004_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3005_ (.D(_0005_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3006_ (.D(_0006_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3007_ (.D(_0032_),
    .CLK(net73),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3008_ (.D(_0033_),
    .CLK(net82),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3009_ (.D(_0034_),
    .CLK(net71),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3010_ (.D(_0035_),
    .CLK(net72),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3011_ (.D(_0036_),
    .CLK(net72),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3012_ (.D(_0037_),
    .CLK(net82),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3013_ (.D(_0038_),
    .CLK(net82),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3014_ (.D(_0039_),
    .CLK(net83),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3015_ (.D(_0040_),
    .CLK(net72),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3016_ (.D(_0041_),
    .CLK(net68),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3017_ (.D(_0042_),
    .CLK(net73),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3018_ (.D(_0043_),
    .CLK(net83),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3019_ (.D(_0044_),
    .CLK(net72),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3020_ (.D(_0045_),
    .CLK(net104),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3021_ (.D(_0046_),
    .CLK(net105),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3022_ (.D(_0047_),
    .CLK(net109),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3023_ (.D(_0048_),
    .CLK(net105),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3024_ (.D(_0049_),
    .CLK(net104),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3025_ (.D(_0050_),
    .CLK(net104),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3026_ (.D(_0051_),
    .CLK(net104),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3027_ (.D(_0052_),
    .CLK(net95),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3028_ (.D(_0053_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3029_ (.D(_0054_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3030_ (.D(_0055_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3031_ (.D(_0056_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3032_ (.D(_0057_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3033_ (.D(_0058_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3034_ (.D(_0059_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3035_ (.D(_0060_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3036_ (.D(_0061_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3037_ (.D(_0062_),
    .CLK(net92),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3038_ (.D(_0063_),
    .CLK(net102),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3039_ (.D(_0064_),
    .CLK(net102),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3040_ (.D(_0065_),
    .CLK(net102),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3041_ (.D(_0066_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3042_ (.D(_0067_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3043_ (.D(_0068_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3044_ (.D(_0069_),
    .CLK(net97),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3045_ (.D(_0070_),
    .CLK(net96),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3046_ (.D(_0071_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3047_ (.D(_0072_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3048_ (.D(_0073_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3049_ (.D(_0074_),
    .CLK(net106),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3050_ (.D(_0075_),
    .CLK(net107),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3051_ (.D(_0076_),
    .CLK(net107),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3052_ (.D(_0077_),
    .CLK(net76),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3053_ (.D(_0078_),
    .CLK(net77),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3054_ (.D(_0079_),
    .CLK(net62),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3055_ (.D(_0080_),
    .CLK(net76),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3056_ (.D(_0081_),
    .CLK(net76),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3057_ (.D(_0082_),
    .CLK(net68),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3058_ (.D(_0083_),
    .CLK(net68),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3059_ (.D(_0084_),
    .CLK(net68),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3060_ (.D(_0085_),
    .CLK(net56),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3061_ (.D(_0086_),
    .CLK(net75),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3062_ (.D(_0087_),
    .CLK(net56),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3063_ (.D(_0088_),
    .CLK(net78),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3064_ (.D(_0089_),
    .CLK(net58),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3065_ (.D(_0090_),
    .CLK(net58),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3066_ (.D(_0091_),
    .CLK(net49),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3067_ (.D(_0092_),
    .CLK(net49),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3068_ (.D(_0093_),
    .CLK(net62),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3069_ (.D(_0094_),
    .CLK(net76),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3070_ (.D(_0095_),
    .CLK(net78),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3071_ (.D(_0096_),
    .CLK(net78),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3072_ (.D(_0097_),
    .CLK(net76),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3073_ (.D(_0098_),
    .CLK(net78),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3074_ (.D(_0099_),
    .CLK(net77),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3075_ (.D(_0100_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3076_ (.D(_0101_),
    .CLK(net56),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3077_ (.D(_0102_),
    .CLK(net57),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3078_ (.D(_0103_),
    .CLK(net57),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3079_ (.D(_0104_),
    .CLK(net58),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3080_ (.D(_0105_),
    .CLK(net58),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3081_ (.D(_0106_),
    .CLK(net47),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3082_ (.D(_0107_),
    .CLK(net48),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3083_ (.D(_0108_),
    .CLK(net48),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3084_ (.D(_0109_),
    .CLK(net62),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3085_ (.D(_0110_),
    .CLK(net78),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3086_ (.D(_0111_),
    .CLK(net69),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3087_ (.D(_0112_),
    .CLK(net67),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3088_ (.D(_0113_),
    .CLK(net109),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3089_ (.D(_0114_),
    .CLK(net110),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3090_ (.D(_0115_),
    .CLK(net110),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3091_ (.D(_0116_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3092_ (.D(_0117_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3093_ (.D(_0118_),
    .CLK(net111),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3094_ (.D(_0119_),
    .CLK(net111),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3095_ (.D(_0120_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3096_ (.D(_0121_),
    .CLK(net115),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3097_ (.D(_0122_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3098_ (.D(_0123_),
    .CLK(net99),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3099_ (.D(_0124_),
    .CLK(net100),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3100_ (.D(_0125_),
    .CLK(net100),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3101_ (.D(_0126_),
    .CLK(net101),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3102_ (.D(_0127_),
    .CLK(net101),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3103_ (.D(_0128_),
    .CLK(net118),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3104_ (.D(_0129_),
    .CLK(net118),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3105_ (.D(_0130_),
    .CLK(net118),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3106_ (.D(_0131_),
    .CLK(net118),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3107_ (.D(_0132_),
    .CLK(net119),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3108_ (.D(_0133_),
    .CLK(net124),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3109_ (.D(_0134_),
    .CLK(net124),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3110_ (.D(_0135_),
    .CLK(net124),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3111_ (.D(_0136_),
    .CLK(net124),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3112_ (.D(_0137_),
    .CLK(net124),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3113_ (.D(_0138_),
    .CLK(net121),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3114_ (.D(_0139_),
    .CLK(net122),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3115_ (.D(_0140_),
    .CLK(net112),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3116_ (.D(_0141_),
    .CLK(net85),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3117_ (.D(_0142_),
    .CLK(net84),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3118_ (.D(_0014_),
    .CLK(net77),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3119_ (.D(_0143_),
    .CLK(net80),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3120_ (.D(_0144_),
    .CLK(net80),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3121_ (.D(_0016_),
    .CLK(net82),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3122_ (.D(_0015_),
    .CLK(net82),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3123_ (.D(_0145_),
    .CLK(net84),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3124_ (.D(_0146_),
    .CLK(net84),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3125_ (.D(_0147_),
    .CLK(net109),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3126_ (.D(_0148_),
    .CLK(net109),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3127_ (.D(_0149_),
    .CLK(net109),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3128_ (.D(_0150_),
    .CLK(net111),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3129_ (.D(_0151_),
    .CLK(net111),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3130_ (.D(_0152_),
    .CLK(net111),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3131_ (.D(_0153_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3132_ (.D(_0154_),
    .CLK(net107),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3133_ (.D(_0155_),
    .CLK(net117),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3134_ (.D(_0156_),
    .CLK(net115),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3135_ (.D(_0157_),
    .CLK(net115),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3136_ (.D(_0158_),
    .CLK(net115),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3137_ (.D(_0159_),
    .CLK(net116),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3138_ (.D(_0160_),
    .CLK(net116),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3139_ (.D(_0161_),
    .CLK(net101),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3140_ (.D(_0162_),
    .CLK(net102),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3141_ (.D(_0163_),
    .CLK(net118),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3142_ (.D(_0164_),
    .CLK(net119),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3143_ (.D(_0165_),
    .CLK(net123),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3144_ (.D(_0166_),
    .CLK(net123),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3145_ (.D(_0167_),
    .CLK(net123),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3146_ (.D(_0168_),
    .CLK(net123),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3147_ (.D(_0169_),
    .CLK(net123),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3148_ (.D(_0170_),
    .CLK(net121),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3149_ (.D(_0171_),
    .CLK(net121),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3150_ (.D(_0172_),
    .CLK(net122),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3151_ (.D(_0173_),
    .CLK(net121),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3152_ (.D(_0174_),
    .CLK(net121),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3153_ (.D(_0175_),
    .CLK(net112),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3154_ (.D(_0176_),
    .CLK(net84),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3155_ (.D(_0013_),
    .CLK(net67),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3156_ (.D(_0177_),
    .CLK(net58),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3157_ (.D(_0178_),
    .CLK(net63),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3158_ (.D(_0179_),
    .CLK(net62),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3159_ (.D(_0180_),
    .CLK(net62),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3160_ (.D(_0181_),
    .CLK(net49),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3161_ (.D(_0182_),
    .CLK(net80),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3162_ (.D(_0183_),
    .CLK(net85),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3163_ (.D(_0184_),
    .CLK(net90),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3164_ (.D(_0185_),
    .CLK(net90),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3165_ (.D(_0186_),
    .CLK(net90),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3166_ (.D(_0187_),
    .CLK(net90),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3167_ (.D(_0188_),
    .CLK(net91),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3168_ (.D(_0189_),
    .CLK(net91),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3169_ (.D(_0190_),
    .CLK(net93),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3170_ (.D(_0191_),
    .CLK(net93),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3171_ (.D(_0192_),
    .CLK(net95),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3172_ (.D(_0193_),
    .CLK(net95),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3173_ (.D(_0194_),
    .CLK(net104),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3174_ (.D(_0195_),
    .CLK(net95),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3175_ (.D(_0196_),
    .CLK(net95),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3176_ (.D(_0197_),
    .CLK(net79),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3177_ (.D(_0198_),
    .CLK(net97),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3178_ (.D(_0199_),
    .CLK(net79),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3179_ (.D(_0200_),
    .CLK(net69),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3180_ (.D(_0201_),
    .CLK(net69),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3181_ (.D(_0202_),
    .CLK(net67),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3182_ (.D(_0203_),
    .CLK(net69),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3183_ (.D(_0204_),
    .CLK(net69),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3184_ (.D(_0205_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3185_ (.D(_0206_),
    .CLK(net71),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3186_ (.D(_0207_),
    .CLK(net70),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3187_ (.D(_0208_),
    .CLK(net77),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3188_ (.D(_0209_),
    .CLK(net71),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3189_ (.D(_0017_),
    .CLK(net54),
    .Q(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3190_ (.D(_0018_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3191_ (.D(_0019_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3192_ (.D(_0020_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3193_ (.D(_0021_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3194_ (.D(_0022_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3195_ (.D(_0023_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3196_ (.D(_0024_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3197_ (.D(_0025_),
    .CLK(net50),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3198_ (.D(_0210_),
    .CLK(net84),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3199_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3200_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3201_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3202_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(net41),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3203_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(net44),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3204_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3205_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3206_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(net52),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3207_ (.D(_0211_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3208_ (.D(_0212_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3209_ (.D(_0213_),
    .CLK(net71),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3210_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(net52),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3211_ (.D(_0214_),
    .CLK(net66),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3212_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3213_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(net40),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3214_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(net41),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3215_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(net43),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3216_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(net44),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3217_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3218_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(net47),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3219_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(net56),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3220_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(net54),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3221_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(net56),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__C (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__B (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__B (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A2 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__B (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__B (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__B2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A2 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A2 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A4 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A3 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__C (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__B (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__B (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__B2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__I (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A3 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__B (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A2 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A2 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__B (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__B (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__B (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A3 (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__B (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__D (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_GWEN  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__D (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A2 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__D (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__D (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__B (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__B (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__B (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A3 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A3 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__B2 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__B (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__C (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__B (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__I (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__I (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__I (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__B (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__I (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__I (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__I (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__S (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_0_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3379_ (.I(\u_scanchain_local.clk_out ),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3380_ (.I(\u_scanchain_local.data_out ),
    .Z(net7));
 gf180mcu_fd_ip_sram__sram256x8m8wm1 \u_cpu.rf_ram.RAM0  (.CEN(net156),
    .CLK(net90),
    .GWEN(_0026_),
    .A({\u_cpu.rf_ram.addr[7] ,
    \u_cpu.rf_ram.addr[6] ,
    \u_cpu.rf_ram.addr[5] ,
    \u_cpu.rf_ram.addr[4] ,
    \u_cpu.rf_ram.addr[3] ,
    \u_cpu.rf_ram.addr[2] ,
    \u_cpu.rf_ram.addr[1] ,
    \u_cpu.rf_ram.addr[0] }),
    .D({\u_cpu.rf_ram.i_wdata[7] ,
    \u_cpu.rf_ram.i_wdata[6] ,
    \u_cpu.rf_ram.i_wdata[5] ,
    \u_cpu.rf_ram.i_wdata[4] ,
    \u_cpu.rf_ram.i_wdata[3] ,
    \u_cpu.rf_ram.i_wdata[2] ,
    \u_cpu.rf_ram.i_wdata[1] ,
    \u_cpu.rf_ram.i_wdata[0] }),
    .Q({\u_cpu.rf_ram.data[7] ,
    \u_cpu.rf_ram.data[6] ,
    \u_cpu.rf_ram.data[5] ,
    \u_cpu.rf_ram.data[4] ,
    \u_cpu.rf_ram.data[3] ,
    \u_cpu.rf_ram.data[2] ,
    \u_cpu.rf_ram.data[1] ,
    \u_cpu.rf_ram.data[0] }),
    .WEN({net11,
    net11,
    net11,
    net11,
    net10,
    net9,
    net9,
    net8}));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.input_buf_clk  (.I(net1),
    .Z(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 \u_scanchain_local.out_flop  (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(net31),
    .Q(\u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.output_buffers[2]  (.I(\u_scanchain_local.data_out_i ),
    .Z(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.output_buffers[3]  (.I(net23),
    .Z(\u_scanchain_local.clk_out ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[0]  (.D(net3),
    .SE(net143),
    .SI(\u_arbiter.o_wb_cpu_cyc ),
    .CLK(net25),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[10]  (.D(\u_arbiter.i_wb_cpu_rdt[7] ),
    .SE(net139),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(net22),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[11]  (.D(\u_arbiter.i_wb_cpu_rdt[8] ),
    .SE(net140),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(net22),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[12]  (.D(\u_arbiter.i_wb_cpu_rdt[9] ),
    .SE(net138),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(net20),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[13]  (.D(\u_arbiter.i_wb_cpu_rdt[10] ),
    .SE(net134),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[14]  (.D(\u_arbiter.i_wb_cpu_rdt[11] ),
    .SE(net138),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(net20),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[15]  (.D(\u_arbiter.i_wb_cpu_rdt[12] ),
    .SE(net135),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[16]  (.D(\u_arbiter.i_wb_cpu_rdt[13] ),
    .SE(net134),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[17]  (.D(\u_arbiter.i_wb_cpu_rdt[14] ),
    .SE(net134),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[18]  (.D(\u_arbiter.i_wb_cpu_rdt[15] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[19]  (.D(\u_arbiter.i_wb_cpu_rdt[16] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[1]  (.D(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .SE(net143),
    .SI(\u_arbiter.o_wb_cpu_we ),
    .CLK(net25),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[20]  (.D(\u_arbiter.i_wb_cpu_rdt[17] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[21]  (.D(\u_arbiter.i_wb_cpu_rdt[18] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(net14),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[22]  (.D(\u_arbiter.i_wb_cpu_rdt[19] ),
    .SE(net131),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[23]  (.D(\u_arbiter.i_wb_cpu_rdt[20] ),
    .SE(net133),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[24]  (.D(\u_arbiter.i_wb_cpu_rdt[21] ),
    .SE(net132),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(net14),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[25]  (.D(\u_arbiter.i_wb_cpu_rdt[22] ),
    .SE(net132),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[26]  (.D(\u_arbiter.i_wb_cpu_rdt[23] ),
    .SE(net133),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[27]  (.D(\u_arbiter.i_wb_cpu_rdt[24] ),
    .SE(net134),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[28]  (.D(\u_arbiter.i_wb_cpu_rdt[25] ),
    .SE(net134),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[29]  (.D(\u_arbiter.i_wb_cpu_rdt[26] ),
    .SE(net135),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[2]  (.D(net12),
    .SE(net139),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[0] ),
    .CLK(net21),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[30]  (.D(\u_arbiter.i_wb_cpu_rdt[27] ),
    .SE(net135),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[31]  (.D(\u_arbiter.i_wb_cpu_rdt[28] ),
    .SE(net135),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[32]  (.D(\u_arbiter.i_wb_cpu_rdt[29] ),
    .SE(net148),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(net30),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[33]  (.D(\u_arbiter.i_wb_cpu_rdt[30] ),
    .SE(net148),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(net30),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[34]  (.D(\u_arbiter.i_wb_cpu_rdt[31] ),
    .SE(net148),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[35]  (.D(\u_scanchain_local.module_data_in[34] ),
    .SE(net148),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[36]  (.D(\u_scanchain_local.module_data_in[35] ),
    .SE(net148),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[37]  (.D(\u_scanchain_local.module_data_in[36] ),
    .SE(net142),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[38]  (.D(\u_scanchain_local.module_data_in[37] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[0] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[39]  (.D(\u_scanchain_local.module_data_in[38] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[1] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[3]  (.D(\u_arbiter.i_wb_cpu_rdt[0] ),
    .SE(net139),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[1] ),
    .CLK(net21),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[40]  (.D(\u_scanchain_local.module_data_in[39] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[2] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[41]  (.D(\u_scanchain_local.module_data_in[40] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[3] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[42]  (.D(\u_scanchain_local.module_data_in[41] ),
    .SE(net141),
    .SI(\u_arbiter.o_wb_cpu_adr[4] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[43]  (.D(\u_scanchain_local.module_data_in[42] ),
    .SE(net142),
    .SI(\u_arbiter.o_wb_cpu_adr[5] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[44]  (.D(\u_scanchain_local.module_data_in[43] ),
    .SE(net151),
    .SI(\u_arbiter.o_wb_cpu_adr[6] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[45]  (.D(\u_scanchain_local.module_data_in[44] ),
    .SE(net151),
    .SI(\u_arbiter.o_wb_cpu_adr[7] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[46]  (.D(\u_scanchain_local.module_data_in[45] ),
    .SE(net150),
    .SI(\u_arbiter.o_wb_cpu_adr[8] ),
    .CLK(net34),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[47]  (.D(\u_scanchain_local.module_data_in[46] ),
    .SE(net150),
    .SI(\u_arbiter.o_wb_cpu_adr[9] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[48]  (.D(\u_scanchain_local.module_data_in[47] ),
    .SE(net145),
    .SI(\u_arbiter.o_wb_cpu_adr[10] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[49]  (.D(\u_scanchain_local.module_data_in[48] ),
    .SE(net145),
    .SI(\u_arbiter.o_wb_cpu_adr[11] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[4]  (.D(\u_arbiter.i_wb_cpu_rdt[1] ),
    .SE(net139),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[2] ),
    .CLK(net21),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[50]  (.D(\u_scanchain_local.module_data_in[49] ),
    .SE(net145),
    .SI(\u_arbiter.o_wb_cpu_adr[12] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[51]  (.D(\u_scanchain_local.module_data_in[50] ),
    .SE(net145),
    .SI(\u_arbiter.o_wb_cpu_adr[13] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[52]  (.D(\u_scanchain_local.module_data_in[51] ),
    .SE(net145),
    .SI(\u_arbiter.o_wb_cpu_adr[14] ),
    .CLK(net28),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[53]  (.D(\u_scanchain_local.module_data_in[52] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[15] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[54]  (.D(\u_scanchain_local.module_data_in[53] ),
    .SE(net136),
    .SI(\u_arbiter.o_wb_cpu_adr[16] ),
    .CLK(net18),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[55]  (.D(\u_scanchain_local.module_data_in[54] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[17] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[56]  (.D(\u_scanchain_local.module_data_in[55] ),
    .SE(net147),
    .SI(\u_arbiter.o_wb_cpu_adr[18] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[57]  (.D(\u_scanchain_local.module_data_in[56] ),
    .SE(net146),
    .SI(\u_arbiter.o_wb_cpu_adr[19] ),
    .CLK(net28),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[58]  (.D(\u_scanchain_local.module_data_in[57] ),
    .SE(net146),
    .SI(\u_arbiter.o_wb_cpu_adr[20] ),
    .CLK(net28),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[59]  (.D(\u_scanchain_local.module_data_in[58] ),
    .SE(net150),
    .SI(\u_arbiter.o_wb_cpu_adr[21] ),
    .CLK(net34),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[5]  (.D(\u_arbiter.i_wb_cpu_rdt[2] ),
    .SE(net139),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[3] ),
    .CLK(net21),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[60]  (.D(\u_scanchain_local.module_data_in[59] ),
    .SE(net150),
    .SI(\u_arbiter.o_wb_cpu_adr[22] ),
    .CLK(net34),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[61]  (.D(\u_scanchain_local.module_data_in[60] ),
    .SE(net149),
    .SI(\u_arbiter.o_wb_cpu_adr[23] ),
    .CLK(net33),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[62]  (.D(\u_scanchain_local.module_data_in[61] ),
    .SE(net149),
    .SI(\u_arbiter.o_wb_cpu_adr[24] ),
    .CLK(net33),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[63]  (.D(\u_scanchain_local.module_data_in[62] ),
    .SE(net149),
    .SI(\u_arbiter.o_wb_cpu_adr[25] ),
    .CLK(net33),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[64]  (.D(\u_scanchain_local.module_data_in[63] ),
    .SE(net152),
    .SI(\u_arbiter.o_wb_cpu_adr[26] ),
    .CLK(net34),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[65]  (.D(\u_scanchain_local.module_data_in[64] ),
    .SE(net149),
    .SI(\u_arbiter.o_wb_cpu_adr[27] ),
    .CLK(net33),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[66]  (.D(\u_scanchain_local.module_data_in[65] ),
    .SE(net149),
    .SI(\u_arbiter.o_wb_cpu_adr[28] ),
    .CLK(net33),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[67]  (.D(\u_scanchain_local.module_data_in[66] ),
    .SE(net151),
    .SI(\u_arbiter.o_wb_cpu_adr[29] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[68]  (.D(\u_scanchain_local.module_data_in[67] ),
    .SE(net151),
    .SI(\u_arbiter.o_wb_cpu_adr[30] ),
    .CLK(net32),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[69]  (.D(\u_scanchain_local.module_data_in[68] ),
    .SE(net151),
    .SI(\u_arbiter.o_wb_cpu_adr[31] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[6]  (.D(\u_arbiter.i_wb_cpu_rdt[3] ),
    .SE(net140),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(net21),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[7]  (.D(\u_arbiter.i_wb_cpu_rdt[4] ),
    .SE(net142),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(net22),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[8]  (.D(\u_arbiter.i_wb_cpu_rdt[5] ),
    .SE(net142),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(net24),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[9]  (.D(\u_arbiter.i_wb_cpu_rdt[6] ),
    .SE(net140),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(net22),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout8 (.I(net10),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout9 (.I(net10),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout10 (.I(net11),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout11 (.I(_0026_),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout12 (.I(\u_arbiter.i_wb_cpu_ack ),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout13 (.I(net15),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout14 (.I(net15),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout15 (.I(net19),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout16 (.I(net18),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout17 (.I(net18),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout18 (.I(net19),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout19 (.I(net20),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout20 (.I(net38),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout21 (.I(net26),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout22 (.I(net26),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout23 (.I(net24),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout24 (.I(net25),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout25 (.I(net26),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout26 (.I(net37),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout27 (.I(net29),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout28 (.I(net29),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout29 (.I(net36),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout30 (.I(net36),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout32 (.I(net35),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout33 (.I(net34),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout34 (.I(net35),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout35 (.I(net36),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout36 (.I(net37),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout38 (.I(\u_scanchain_local.clk ),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout39 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net42),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net43),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout44 (.I(net130),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout45 (.I(net50),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net50),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net61),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout51 (.I(net55),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net55),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net55),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net60),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout56 (.I(net59),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net59),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout58 (.I(net60),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net60),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net61),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net64),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout62 (.I(net64),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net89),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net67),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout68 (.I(net75),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout69 (.I(net74),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net74),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout71 (.I(net73),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net74),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net88),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout77 (.I(net81),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout78 (.I(net80),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout79 (.I(net80),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net87),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout82 (.I(net86),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net86),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout84 (.I(net86),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net129),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 fanout90 (.I(net94),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout91 (.I(net94),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout92 (.I(net94),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout94 (.I(net98),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout95 (.I(net97),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net97),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout97 (.I(net98),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout98 (.I(net103),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout99 (.I(net101),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout100 (.I(net101),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout101 (.I(net102),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout102 (.I(net103),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net128),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout104 (.I(net108),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout105 (.I(net108),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net108),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net114),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net113),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout110 (.I(net113),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout114 (.I(net127),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout115 (.I(net117),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout117 (.I(net120),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net120),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net120),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout120 (.I(net126),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout121 (.I(net125),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout122 (.I(net125),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net125),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout124 (.I(net125),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout125 (.I(net126),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net127),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net128),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout128 (.I(net129),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net5),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout131 (.I(net133),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout132 (.I(net133),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout133 (.I(net137),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout134 (.I(net136),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout135 (.I(net136),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout137 (.I(net138),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout138 (.I(net155),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout139 (.I(net144),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout140 (.I(net144),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout142 (.I(net143),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout143 (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net154),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout145 (.I(net147),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net147),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout147 (.I(net153),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout148 (.I(net153),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout150 (.I(net152),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout151 (.I(net153),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout152 (.I(net153),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout153 (.I(net154),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout154 (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout155 (.I(net4),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_cpu.rf_ram.RAM0_156  (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__B (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__B1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__B1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__B1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__B1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__B1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__B (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__C1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__C1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__C (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__B1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__B1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__B1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__B1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__B1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__B1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__C1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__B1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__B1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__B1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__B1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__B1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__C1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__C1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__C1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__C1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__C1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__B1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__B1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__B1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__B1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__B1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__B1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__B1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__B1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__B1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__C (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__C (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__B (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A3 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__S (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A3 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__I (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__B (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__C (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__C (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__B2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__B1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__B1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__I (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__B1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__C (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__I (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__B2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__C (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__B (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__B2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__C (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__I (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__B2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__B1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__B1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__B2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__I (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__C (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__C (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__C (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__C (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__B2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__I (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__I (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__B2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__I (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__B2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__B2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__C (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__B (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__B (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__B (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__C (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__C (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__B1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__B2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__B2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__B (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A3 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A3 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__C (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__B (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__B (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__B (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__B1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__B1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__B2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__B2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__C (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__B2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__B2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__B1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__B1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A3 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__C (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__B2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__C (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__C (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__B (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__B2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A4 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A3 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A3 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__C (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__B (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__B (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__B2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__B1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__B1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__B1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__B1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__B2 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__B2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__B1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__C (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__B (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__C (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__B2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__C (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__B (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__C (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__C (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__B1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__B2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__B (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__B (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__C (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__B (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__B (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__B2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__B (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__B1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__B2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__B (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__C (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__B (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A3 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__C (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__C (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__B (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__C (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__B2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__C (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__B (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__C2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__S (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__S (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__S (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__S (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__S (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__S (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__S (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A3 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__B2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__B (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__B (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__B2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__B2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__B (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__B2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__C (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__C (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__B2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__B2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__C2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__B (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A3 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__C (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__C1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__B (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__B (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__C1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__B1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__B2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__B2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__B2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__B1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__B2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__C1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__B1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__C2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A3 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__B1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__C (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__C (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__B1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__B (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__B (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__B (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__B2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__C (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__C (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A3 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__S (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__S (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__S (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__S (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__S (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__S (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__S (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__S (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__S (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__S (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__S (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__S (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__S (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__B1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__B1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__B1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__B1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__B1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__B1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__B1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A3 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__S (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__S (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__S (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__S (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__S (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__S (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__S (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__B (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__I (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__S1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__I (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A3 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__I (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__I (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__C (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__B1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__B2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A4 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__B1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__B2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1572__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__B2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__C (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__B1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__B1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__B1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__B1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__S (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__S (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__S (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A4 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__A3 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__I (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__S (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__S (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__I (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__S (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__S (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__S (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__I (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__S (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__S (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__S (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__I (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__S (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__B (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__B (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__B (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A4 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A3 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A3 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A3 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A3 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A3 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A3 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A4 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__A3 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A2 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A2 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A3 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A4 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A3 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__B2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A4 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A3 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A3 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__I (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__I (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A3 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__I0 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__I (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__C (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A1 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A3 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A3 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__B (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__S (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__S (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__B (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__B2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__I (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__B2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A3 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A4 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__B2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__B (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A3 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A4 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__B (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__B (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A3 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__C (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__I (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__C (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A1 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__I0 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__B2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A3 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__B (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A4 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__C (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__A3 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A3 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__B1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__B2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__I0 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__B (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__C (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__S (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__S (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__S (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__S (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__S (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A3 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__S (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__S (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__I1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__I1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__S (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__S (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__S (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__S (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__S (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__I1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__I1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__I1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__I1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__I1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__I1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__I (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__I (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__B1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__B1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__B2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout12_I (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__I (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__I (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__I (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__C2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__B (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__I (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__B2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_D  (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_D  (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_D  (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_D  (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__I1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_D  (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_D  (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_D  (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_D  (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_D  (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_D  (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_D  (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A2 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_D  (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__I1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__I0 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A2 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_D  (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_D  (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_D  (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_D  (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_D  (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_D  (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_D  (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_D  (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_D  (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_D  (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A2 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_D  (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__I1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__I0 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_D  (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_D  (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_D  (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A2 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_D  (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_D  (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A2 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_D  (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A2 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_D  (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_D  (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__I1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__C (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__S0 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__I (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__I (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__I (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__I (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A2 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A1 (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__I (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__I (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__S (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A1 (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_D  (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A3 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__I0 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__B2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__I (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A4 (.I(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__I (.I(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A3 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__B2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__B2 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A2 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__B (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__I (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A2 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__I (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__D (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__I1 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__D (.I(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__C (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A2 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__I (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[0]  (.I(\u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[1]  (.I(\u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[2]  (.I(\u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[3]  (.I(\u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[4]  (.I(\u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[5]  (.I(\u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[6]  (.I(\u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_A[7]  (.I(\u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A1 (.I(\u_cpu.rf_ram.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__I1 (.I(\u_cpu.rf_ram.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__I1 (.I(\u_cpu.rf_ram.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__I1 (.I(\u_cpu.rf_ram.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__I1 (.I(\u_cpu.rf_ram.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__I1 (.I(\u_cpu.rf_ram.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__I1 (.I(\u_cpu.rf_ram.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__I1 (.I(\u_cpu.rf_ram.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[0]  (.I(\u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[1]  (.I(\u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[2]  (.I(\u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[3]  (.I(\u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[4]  (.I(\u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[5]  (.I(\u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[6]  (.I(\u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_D[7]  (.I(\u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__B (.I(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__I (.I(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__B (.I(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__S (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__D (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__D (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__D (.I(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__D (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__D (.I(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__D (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__I0 (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_D  (.I(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_D  (.I(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.input_buf_clk_I  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__B (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__S (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__B (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[0]  (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[3]  (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout8_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout9_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[4]  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[5]  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[6]  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_WEN[7]  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout10_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_D  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout13_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout14_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_CLK  (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout16_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout17_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout15_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout19_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.output_buffers[3]_I  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout23_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout24_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_CLK  (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_CLK  (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout27_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_CLK  (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_CLK  (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_CLK  (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_CLK  (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_CLKN  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_CLK  (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_CLK  (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_CLK  (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_CLK  (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_CLK  (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_CLK  (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_CLK  (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_CLK  (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_CLK  (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_CLK  (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout26_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__CLK (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__CLK (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_cpu.rf_ram.RAM0_CLK  (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__CLK (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_SE  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_SE  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_SE  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_SE  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_SE  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SE  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_SE  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_SE  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_SE  (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_SE  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SE  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_SE  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SE  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_SE  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_SE  (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SE  (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_SE  (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_SE  (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_SE  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_SE  (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_SE  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SE  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_SE  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_SE  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_SE  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_SE  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_SE  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_SE  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_SE  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_SE  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_SE  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_SE  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_SE  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_SE  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SE  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_SE  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_SE  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_SE  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_SE  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout151_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1223 ();
 assign io_oeb[0] = net157;
 assign io_oeb[1] = net158;
 assign io_oeb[2] = net159;
 assign io_oeb[3] = net160;
 assign io_oeb[4] = net161;
 assign io_out[2] = net162;
 assign io_out[3] = net163;
 assign io_out[4] = net164;
endmodule

